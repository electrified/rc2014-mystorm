// Reading file 'chip.asc'..

module chip (output io_0_16_0, output io_0_16_1, input io_16_33_1, input io_0_27_1, output io_0_11_1, input io_0_28_0, output io_0_11_0, output io_0_18_1, output io_0_17_1, output io_0_17_0, input io_33_29_1, output io_0_20_0, output io_0_20_1, output io_0_18_0, input io_33_31_0, output io_0_22_0, output io_0_22_1, input io_0_27_0, input io_0_25_0, input io_3_33_1, input io_4_33_0, input io_33_30_1, input io_30_33_1, input io_31_33_0, input io_31_33_1, input io_30_33_0, input io_33_30_0, input io_33_27_1, input io_29_0_0, input io_33_23_1, input io_33_20_1, input io_33_21_1, input io_33_28_0, input io_33_21_0, output io_31_0_1);

wire n1;
// (0, 0, 'glb_netwk_0')
// (16, 1, 'sp4_r_v_b_36')
// (16, 2, 'sp4_r_v_b_25')
// (16, 3, 'sp4_r_v_b_12')
// (16, 4, 'sp4_r_v_b_1')
// (16, 5, 'sp4_r_v_b_36')
// (16, 6, 'sp4_r_v_b_25')
// (16, 7, 'sp4_r_v_b_12')
// (16, 8, 'sp4_r_v_b_1')
// (16, 9, 'sp4_r_v_b_36')
// (16, 10, 'neigh_op_tnr_6')
// (16, 10, 'sp4_r_v_b_25')
// (16, 11, 'lutff_global/s_r')
// (16, 11, 'neigh_op_rgt_6')
// (16, 11, 'sp4_r_v_b_12')
// (16, 12, 'lutff_global/s_r')
// (16, 12, 'neigh_op_bnr_6')
// (16, 12, 'sp4_r_v_b_1')
// (17, 0, 'fabout')
// (17, 0, 'local_g1_4')
// (17, 0, 'span4_vert_36')
// (17, 1, 'sp4_v_b_36')
// (17, 2, 'sp4_v_b_25')
// (17, 3, 'sp4_v_b_12')
// (17, 4, 'sp4_v_b_1')
// (17, 4, 'sp4_v_t_36')
// (17, 5, 'sp4_v_b_36')
// (17, 6, 'sp4_v_b_25')
// (17, 7, 'sp4_v_b_12')
// (17, 8, 'sp4_v_b_1')
// (17, 8, 'sp4_v_t_36')
// (17, 9, 'sp4_v_b_36')
// (17, 10, 'neigh_op_top_6')
// (17, 10, 'sp4_v_b_25')
// (17, 11, 'lutff_6/out')
// (17, 11, 'lutff_global/s_r')
// (17, 11, 'sp4_v_b_12')
// (17, 12, 'local_g1_6')
// (17, 12, 'lutff_3/in_2')
// (17, 12, 'neigh_op_bot_6')
// (17, 12, 'sp4_v_b_1')
// (18, 10, 'local_g2_6')
// (18, 10, 'lutff_7/in_1')
// (18, 10, 'lutff_global/s_r')
// (18, 10, 'neigh_op_tnl_6')
// (18, 11, 'neigh_op_lft_6')
// (18, 12, 'neigh_op_bnl_6')

wire io_0_16_0;
assign io_0_16_1 = io_0_16_0;
// (0, 0, 'glb_netwk_3')
// (0, 16, 'io_0/D_OUT_0')
// (0, 16, 'io_0/PAD')
// (0, 16, 'io_1/D_OUT_0')
// (0, 16, 'io_1/PAD')
// (0, 16, 'local_g0_7')
// (0, 16, 'local_g1_7')
// (0, 16, 'span4_horz_7')
// (0, 16, 'span4_vert_t_13')
// (0, 17, 'fabout')
// (0, 17, 'local_g0_5')
// (0, 17, 'span4_vert_b_13')
// (0, 18, 'span4_vert_b_9')
// (0, 19, 'span4_vert_b_5')
// (0, 20, 'span4_horz_7')
// (0, 20, 'span4_vert_b_1')
// (1, 16, 'sp4_h_r_18')
// (1, 20, 'sp4_h_r_18')
// (2, 16, 'sp4_h_r_31')
// (2, 20, 'sp4_h_r_31')
// (3, 16, 'sp4_h_r_42')
// (3, 20, 'sp4_h_r_42')
// (4, 16, 'sp4_h_l_42')
// (4, 16, 'sp4_h_r_11')
// (4, 20, 'sp4_h_l_42')
// (4, 20, 'sp4_h_r_11')
// (5, 16, 'sp4_h_r_22')
// (5, 20, 'sp4_h_r_22')
// (6, 16, 'sp4_h_r_35')
// (6, 20, 'sp4_h_r_35')
// (7, 16, 'sp4_h_r_46')
// (7, 20, 'sp4_h_r_46')
// (7, 24, 'sp4_r_v_b_43')
// (7, 25, 'sp4_r_v_b_30')
// (7, 25, 'sp4_r_v_b_46')
// (7, 26, 'sp4_r_v_b_19')
// (7, 26, 'sp4_r_v_b_35')
// (7, 27, 'sp4_r_v_b_22')
// (7, 27, 'sp4_r_v_b_6')
// (7, 28, 'sp4_r_v_b_11')
// (8, 11, 'sp12_v_t_23')
// (8, 12, 'sp12_v_b_23')
// (8, 13, 'sp12_v_b_20')
// (8, 14, 'sp12_v_b_19')
// (8, 15, 'sp12_v_b_16')
// (8, 16, 'local_g1_3')
// (8, 16, 'ram/WCLK')
// (8, 16, 'ram/WCLKE')
// (8, 16, 'sp12_v_b_15')
// (8, 16, 'sp4_h_l_46')
// (8, 16, 'sp4_h_r_11')
// (8, 16, 'sp4_r_v_b_43')
// (8, 17, 'sp12_v_b_12')
// (8, 17, 'sp4_r_v_b_30')
// (8, 18, 'local_g3_3')
// (8, 18, 'ram/WCLK')
// (8, 18, 'ram/WCLKE')
// (8, 18, 'sp12_v_b_11')
// (8, 18, 'sp4_r_v_b_19')
// (8, 19, 'sp12_v_b_8')
// (8, 19, 'sp4_r_v_b_6')
// (8, 20, 'local_g1_3')
// (8, 20, 'ram/WCLK')
// (8, 20, 'ram/WCLKE')
// (8, 20, 'sp12_v_b_7')
// (8, 20, 'sp4_h_l_46')
// (8, 20, 'sp4_h_r_11')
// (8, 21, 'sp12_v_b_4')
// (8, 22, 'local_g3_3')
// (8, 22, 'ram/WCLK')
// (8, 22, 'ram/WCLKE')
// (8, 22, 'sp12_v_b_3')
// (8, 23, 'sp12_h_r_0')
// (8, 23, 'sp12_v_b_0')
// (8, 23, 'sp12_v_t_23')
// (8, 23, 'sp4_h_r_0')
// (8, 23, 'sp4_v_t_43')
// (8, 24, 'local_g0_2')
// (8, 24, 'ram/WCLK')
// (8, 24, 'ram/WCLKE')
// (8, 24, 'sp12_v_b_23')
// (8, 24, 'sp4_h_r_10')
// (8, 24, 'sp4_h_r_5')
// (8, 24, 'sp4_v_b_43')
// (8, 24, 'sp4_v_t_46')
// (8, 25, 'sp12_v_b_20')
// (8, 25, 'sp4_v_b_30')
// (8, 25, 'sp4_v_b_46')
// (8, 26, 'local_g1_3')
// (8, 26, 'ram/WCLK')
// (8, 26, 'ram/WCLKE')
// (8, 26, 'sp12_v_b_19')
// (8, 26, 'sp4_v_b_19')
// (8, 26, 'sp4_v_b_35')
// (8, 27, 'sp12_v_b_16')
// (8, 27, 'sp4_v_b_22')
// (8, 27, 'sp4_v_b_6')
// (8, 28, 'local_g1_3')
// (8, 28, 'ram/WCLK')
// (8, 28, 'ram/WCLKE')
// (8, 28, 'sp12_v_b_15')
// (8, 28, 'sp4_v_b_11')
// (8, 29, 'sp12_v_b_12')
// (8, 30, 'local_g3_3')
// (8, 30, 'ram/WCLK')
// (8, 30, 'ram/WCLKE')
// (8, 30, 'sp12_v_b_11')
// (8, 31, 'sp12_v_b_8')
// (8, 32, 'sp12_v_b_7')
// (8, 33, 'span12_vert_4')
// (9, 15, 'sp4_v_t_43')
// (9, 16, 'sp4_h_r_22')
// (9, 16, 'sp4_v_b_43')
// (9, 17, 'sp4_v_b_30')
// (9, 18, 'sp4_v_b_19')
// (9, 19, 'sp4_h_r_1')
// (9, 19, 'sp4_v_b_6')
// (9, 20, 'sp4_h_r_22')
// (9, 23, 'sp12_h_r_3')
// (9, 23, 'sp4_h_r_13')
// (9, 24, 'sp4_h_r_16')
// (9, 24, 'sp4_h_r_23')
// (10, 16, 'sp4_h_r_35')
// (10, 19, 'sp4_h_r_12')
// (10, 20, 'sp4_h_r_35')
// (10, 23, 'sp12_h_r_4')
// (10, 23, 'sp4_h_r_24')
// (10, 23, 'sp4_h_r_8')
// (10, 24, 'sp4_h_r_29')
// (10, 24, 'sp4_h_r_34')
// (11, 16, 'sp4_h_r_46')
// (11, 17, 'sp4_r_v_b_40')
// (11, 18, 'sp4_r_v_b_29')
// (11, 19, 'sp4_h_r_25')
// (11, 19, 'sp4_r_v_b_16')
// (11, 20, 'sp4_h_r_46')
// (11, 20, 'sp4_r_v_b_5')
// (11, 21, 'sp4_r_v_b_40')
// (11, 22, 'neigh_op_tnr_0')
// (11, 22, 'sp4_r_v_b_29')
// (11, 23, 'neigh_op_rgt_0')
// (11, 23, 'sp12_h_r_7')
// (11, 23, 'sp4_h_r_21')
// (11, 23, 'sp4_h_r_37')
// (11, 23, 'sp4_r_v_b_16')
// (11, 24, 'neigh_op_bnr_0')
// (11, 24, 'sp4_h_r_40')
// (11, 24, 'sp4_h_r_47')
// (11, 24, 'sp4_r_v_b_5')
// (12, 16, 'sp4_h_l_46')
// (12, 16, 'sp4_v_t_40')
// (12, 17, 'sp4_v_b_40')
// (12, 18, 'sp4_v_b_29')
// (12, 19, 'sp4_h_r_36')
// (12, 19, 'sp4_v_b_16')
// (12, 20, 'sp4_h_l_46')
// (12, 20, 'sp4_r_v_b_36')
// (12, 20, 'sp4_v_b_5')
// (12, 20, 'sp4_v_t_40')
// (12, 21, 'sp4_r_v_b_25')
// (12, 21, 'sp4_r_v_b_41')
// (12, 21, 'sp4_v_b_40')
// (12, 22, 'neigh_op_top_0')
// (12, 22, 'sp4_r_v_b_12')
// (12, 22, 'sp4_r_v_b_28')
// (12, 22, 'sp4_v_b_29')
// (12, 23, 'lutff_0/out')
// (12, 23, 'sp12_h_r_8')
// (12, 23, 'sp4_h_l_37')
// (12, 23, 'sp4_h_r_0')
// (12, 23, 'sp4_h_r_32')
// (12, 23, 'sp4_r_v_b_1')
// (12, 23, 'sp4_r_v_b_17')
// (12, 23, 'sp4_v_b_16')
// (12, 24, 'neigh_op_bot_0')
// (12, 24, 'sp4_h_l_40')
// (12, 24, 'sp4_h_l_47')
// (12, 24, 'sp4_r_v_b_4')
// (12, 24, 'sp4_v_b_5')
// (13, 19, 'sp4_h_l_36')
// (13, 19, 'sp4_h_r_1')
// (13, 19, 'sp4_v_t_36')
// (13, 20, 'sp4_h_r_9')
// (13, 20, 'sp4_v_b_36')
// (13, 20, 'sp4_v_t_41')
// (13, 21, 'sp4_v_b_25')
// (13, 21, 'sp4_v_b_41')
// (13, 22, 'neigh_op_tnl_0')
// (13, 22, 'sp4_v_b_12')
// (13, 22, 'sp4_v_b_28')
// (13, 23, 'neigh_op_lft_0')
// (13, 23, 'sp12_h_r_11')
// (13, 23, 'sp4_h_r_13')
// (13, 23, 'sp4_h_r_45')
// (13, 23, 'sp4_v_b_1')
// (13, 23, 'sp4_v_b_17')
// (13, 24, 'neigh_op_bnl_0')
// (13, 24, 'sp4_h_r_10')
// (13, 24, 'sp4_v_b_4')
// (14, 19, 'sp4_h_r_12')
// (14, 20, 'sp4_h_r_20')
// (14, 23, 'sp12_h_r_12')
// (14, 23, 'sp4_h_l_45')
// (14, 23, 'sp4_h_r_11')
// (14, 23, 'sp4_h_r_24')
// (14, 24, 'sp4_h_r_23')
// (15, 19, 'sp4_h_r_25')
// (15, 20, 'sp4_h_r_33')
// (15, 23, 'sp12_h_r_15')
// (15, 23, 'sp4_h_r_22')
// (15, 23, 'sp4_h_r_37')
// (15, 24, 'sp4_h_r_34')
// (16, 19, 'sp4_h_r_36')
// (16, 20, 'sp4_h_r_44')
// (16, 23, 'sp12_h_r_16')
// (16, 23, 'sp4_h_l_37')
// (16, 23, 'sp4_h_r_35')
// (16, 24, 'sp4_h_r_47')
// (17, 19, 'sp4_h_l_36')
// (17, 19, 'sp4_h_r_4')
// (17, 20, 'sp4_h_l_44')
// (17, 20, 'sp4_h_r_0')
// (17, 23, 'sp12_h_r_19')
// (17, 23, 'sp4_h_r_46')
// (17, 24, 'sp4_h_l_47')
// (17, 24, 'sp4_h_r_10')
// (18, 19, 'sp4_h_r_17')
// (18, 20, 'sp4_h_r_13')
// (18, 23, 'sp12_h_r_20')
// (18, 23, 'sp4_h_l_46')
// (18, 23, 'sp4_h_r_2')
// (18, 24, 'sp4_h_r_23')
// (19, 19, 'sp4_h_r_28')
// (19, 20, 'sp4_h_r_24')
// (19, 23, 'sp12_h_r_23')
// (19, 23, 'sp4_h_r_15')
// (19, 24, 'sp4_h_r_34')
// (20, 19, 'sp4_h_r_41')
// (20, 20, 'sp4_h_r_37')
// (20, 23, 'sp12_h_l_23')
// (20, 23, 'sp4_h_r_26')
// (20, 24, 'sp4_h_r_47')
// (21, 19, 'sp4_h_l_41')
// (21, 19, 'sp4_h_r_0')
// (21, 20, 'sp4_h_l_37')
// (21, 20, 'sp4_h_r_8')
// (21, 23, 'sp4_h_r_39')
// (21, 24, 'sp4_h_l_47')
// (21, 24, 'sp4_h_r_10')
// (22, 19, 'sp4_h_r_13')
// (22, 20, 'sp4_h_r_21')
// (22, 23, 'sp4_h_l_39')
// (22, 23, 'sp4_h_r_10')
// (22, 24, 'sp4_h_r_23')
// (23, 19, 'sp4_h_r_24')
// (23, 20, 'sp4_h_r_32')
// (23, 23, 'sp4_h_r_23')
// (23, 24, 'sp4_h_r_34')
// (24, 16, 'sp4_r_v_b_43')
// (24, 17, 'sp4_r_v_b_30')
// (24, 18, 'sp4_r_v_b_19')
// (24, 19, 'sp4_h_r_37')
// (24, 19, 'sp4_r_v_b_6')
// (24, 20, 'sp4_h_r_45')
// (24, 23, 'sp4_h_r_34')
// (24, 24, 'sp4_h_r_47')
// (25, 15, 'sp4_v_t_43')
// (25, 16, 'local_g3_3')
// (25, 16, 'ram/WCLK')
// (25, 16, 'ram/WCLKE')
// (25, 16, 'sp4_v_b_43')
// (25, 17, 'sp4_v_b_30')
// (25, 18, 'local_g1_3')
// (25, 18, 'ram/WCLK')
// (25, 18, 'ram/WCLKE')
// (25, 18, 'sp4_v_b_19')
// (25, 19, 'sp4_h_l_37')
// (25, 19, 'sp4_v_b_6')
// (25, 20, 'local_g1_3')
// (25, 20, 'ram/WCLK')
// (25, 20, 'ram/WCLKE')
// (25, 20, 'sp4_h_l_45')
// (25, 20, 'sp4_h_r_11')
// (25, 20, 'sp4_r_v_b_43')
// (25, 21, 'sp4_r_v_b_30')
// (25, 22, 'local_g3_3')
// (25, 22, 'ram/WCLK')
// (25, 22, 'ram/WCLKE')
// (25, 22, 'sp4_r_v_b_19')
// (25, 23, 'sp4_h_r_47')
// (25, 23, 'sp4_r_v_b_6')
// (25, 24, 'local_g0_2')
// (25, 24, 'ram/WCLK')
// (25, 24, 'ram/WCLKE')
// (25, 24, 'sp4_h_l_47')
// (25, 24, 'sp4_h_r_10')
// (25, 24, 'sp4_r_v_b_38')
// (25, 24, 'sp4_r_v_b_43')
// (25, 25, 'sp4_r_v_b_27')
// (25, 25, 'sp4_r_v_b_30')
// (25, 26, 'local_g3_3')
// (25, 26, 'ram/WCLK')
// (25, 26, 'ram/WCLKE')
// (25, 26, 'sp4_r_v_b_14')
// (25, 26, 'sp4_r_v_b_19')
// (25, 27, 'sp4_r_v_b_3')
// (25, 27, 'sp4_r_v_b_6')
// (25, 28, 'local_g3_3')
// (25, 28, 'ram/WCLK')
// (25, 28, 'ram/WCLKE')
// (25, 28, 'sp4_r_v_b_43')
// (25, 29, 'sp4_r_v_b_30')
// (25, 30, 'local_g3_3')
// (25, 30, 'ram/WCLK')
// (25, 30, 'ram/WCLKE')
// (25, 30, 'sp4_r_v_b_19')
// (25, 31, 'sp4_r_v_b_6')
// (26, 19, 'sp4_v_t_43')
// (26, 20, 'sp4_h_r_22')
// (26, 20, 'sp4_v_b_43')
// (26, 21, 'sp4_v_b_30')
// (26, 22, 'sp4_v_b_19')
// (26, 23, 'sp4_h_l_47')
// (26, 23, 'sp4_h_r_6')
// (26, 23, 'sp4_v_b_6')
// (26, 23, 'sp4_v_t_38')
// (26, 23, 'sp4_v_t_43')
// (26, 24, 'sp4_h_r_23')
// (26, 24, 'sp4_v_b_38')
// (26, 24, 'sp4_v_b_43')
// (26, 25, 'sp4_v_b_27')
// (26, 25, 'sp4_v_b_30')
// (26, 26, 'sp4_v_b_14')
// (26, 26, 'sp4_v_b_19')
// (26, 27, 'sp4_v_b_3')
// (26, 27, 'sp4_v_b_6')
// (26, 27, 'sp4_v_t_43')
// (26, 28, 'sp4_v_b_43')
// (26, 29, 'sp4_v_b_30')
// (26, 30, 'sp4_v_b_19')
// (26, 31, 'sp4_v_b_6')
// (27, 20, 'sp4_h_r_35')
// (27, 23, 'sp4_h_r_19')
// (27, 24, 'sp4_h_r_34')
// (28, 20, 'sp4_h_r_46')
// (28, 23, 'sp4_h_r_30')
// (28, 24, 'sp4_h_r_47')
// (29, 20, 'sp4_h_l_46')
// (29, 23, 'sp4_h_r_43')
// (29, 24, 'sp4_h_l_47')
// (30, 23, 'sp4_h_l_43')

wire io_16_33_1;
// (0, 0, 'glb_netwk_4')
// (15, 15, 'lutff_global/clk')
// (15, 32, 'neigh_op_tnr_2')
// (15, 32, 'neigh_op_tnr_6')
// (16, 13, 'lutff_global/clk')
// (16, 14, 'lutff_global/clk')
// (16, 15, 'lutff_global/clk')
// (16, 32, 'neigh_op_top_2')
// (16, 32, 'neigh_op_top_6')
// (16, 33, 'fabout')
// (16, 33, 'io_1/D_IN_0')
// (16, 33, 'io_1/PAD')
// (16, 33, 'local_g1_2')
// (16, 33, 'span4_horz_r_2')
// (17, 32, 'neigh_op_tnl_2')
// (17, 32, 'neigh_op_tnl_6')
// (17, 33, 'span4_horz_r_6')
// (18, 33, 'span4_horz_r_10')
// (19, 33, 'span4_horz_r_14')
// (20, 33, 'span4_horz_l_14')

reg n4 = 0;
// (0, 0, 'glb_netwk_5')
// (6, 20, 'lutff_global/clk')
// (6, 21, 'lutff_global/clk')
// (7, 19, 'lutff_global/clk')
// (7, 20, 'lutff_global/clk')
// (7, 21, 'lutff_global/clk')
// (7, 22, 'lutff_global/clk')
// (15, 1, 'sp4_r_v_b_9')
// (15, 2, 'sp4_r_v_b_43')
// (15, 3, 'sp4_r_v_b_30')
// (15, 4, 'sp4_r_v_b_19')
// (15, 5, 'sp4_r_v_b_6')
// (15, 6, 'sp4_r_v_b_47')
// (15, 7, 'sp4_r_v_b_34')
// (15, 8, 'sp4_r_v_b_23')
// (15, 9, 'sp4_r_v_b_10')
// (15, 10, 'sp4_r_v_b_47')
// (15, 11, 'sp4_r_v_b_34')
// (15, 12, 'neigh_op_tnr_5')
// (15, 12, 'sp4_r_v_b_23')
// (15, 13, 'neigh_op_rgt_5')
// (15, 13, 'sp4_r_v_b_10')
// (15, 14, 'neigh_op_bnr_5')
// (16, 0, 'fabout')
// (16, 0, 'local_g0_1')
// (16, 0, 'span4_vert_9')
// (16, 1, 'sp4_v_b_9')
// (16, 1, 'sp4_v_t_43')
// (16, 2, 'sp4_v_b_43')
// (16, 3, 'sp4_v_b_30')
// (16, 4, 'sp4_v_b_19')
// (16, 5, 'sp4_v_b_6')
// (16, 5, 'sp4_v_t_47')
// (16, 6, 'sp4_v_b_47')
// (16, 7, 'sp4_v_b_34')
// (16, 8, 'sp4_v_b_23')
// (16, 9, 'sp4_v_b_10')
// (16, 9, 'sp4_v_t_47')
// (16, 10, 'sp4_v_b_47')
// (16, 11, 'lutff_global/clk')
// (16, 11, 'sp4_v_b_34')
// (16, 12, 'lutff_global/clk')
// (16, 12, 'neigh_op_top_5')
// (16, 12, 'sp4_v_b_23')
// (16, 13, 'local_g0_5')
// (16, 13, 'lutff_5/in_0')
// (16, 13, 'lutff_5/out')
// (16, 13, 'sp4_v_b_10')
// (16, 14, 'local_g1_5')
// (16, 14, 'lutff_4/in_0')
// (16, 14, 'neigh_op_bot_5')
// (17, 11, 'lutff_global/clk')
// (17, 12, 'neigh_op_tnl_5')
// (17, 13, 'neigh_op_lft_5')
// (17, 14, 'neigh_op_bnl_5')
// (18, 10, 'lutff_global/clk')

wire io_0_27_1;
// (0, 0, 'glb_netwk_6')
// (0, 15, 'span4_vert_t_14')
// (0, 16, 'fabout')
// (0, 16, 'local_g1_6')
// (0, 16, 'span4_vert_b_14')
// (0, 17, 'span4_vert_b_10')
// (0, 18, 'span4_vert_b_6')
// (0, 19, 'span4_vert_b_2')
// (0, 19, 'span4_vert_t_14')
// (0, 20, 'span4_vert_b_14')
// (0, 21, 'span4_vert_b_10')
// (0, 22, 'span4_vert_b_6')
// (0, 23, 'span4_vert_b_2')
// (0, 23, 'span4_vert_t_14')
// (0, 24, 'span4_vert_b_14')
// (0, 25, 'span4_vert_b_10')
// (0, 26, 'span4_vert_b_6')
// (0, 27, 'io_1/D_IN_0')
// (0, 27, 'io_1/PAD')
// (0, 27, 'span12_horz_4')
// (0, 27, 'span4_vert_b_2')
// (1, 26, 'neigh_op_tnl_2')
// (1, 26, 'neigh_op_tnl_6')
// (1, 27, 'neigh_op_lft_2')
// (1, 27, 'neigh_op_lft_6')
// (1, 27, 'sp12_h_r_7')
// (1, 28, 'neigh_op_bnl_2')
// (1, 28, 'neigh_op_bnl_6')
// (2, 27, 'sp12_h_r_8')
// (3, 27, 'sp12_h_r_11')
// (4, 27, 'sp12_h_r_12')
// (5, 27, 'sp12_h_r_15')
// (6, 27, 'sp12_h_r_16')
// (7, 27, 'sp12_h_r_19')
// (8, 15, 'ram/RCLK')
// (8, 17, 'ram/RCLK')
// (8, 19, 'ram/RCLK')
// (8, 21, 'ram/RCLK')
// (8, 23, 'ram/RCLK')
// (8, 25, 'ram/RCLK')
// (8, 27, 'ram/RCLK')
// (8, 27, 'sp12_h_r_20')
// (8, 29, 'ram/RCLK')
// (9, 16, 'sp4_r_v_b_45')
// (9, 17, 'sp4_r_v_b_32')
// (9, 18, 'sp4_r_v_b_21')
// (9, 19, 'sp4_r_v_b_8')
// (9, 27, 'sp12_h_r_23')
// (10, 15, 'sp12_v_t_23')
// (10, 15, 'sp4_h_r_8')
// (10, 15, 'sp4_v_t_45')
// (10, 16, 'sp12_v_b_23')
// (10, 16, 'sp4_v_b_45')
// (10, 17, 'sp12_v_b_20')
// (10, 17, 'sp4_v_b_32')
// (10, 18, 'sp12_v_b_19')
// (10, 18, 'sp4_v_b_21')
// (10, 19, 'sp12_v_b_16')
// (10, 19, 'sp4_v_b_8')
// (10, 20, 'sp12_v_b_15')
// (10, 21, 'sp12_v_b_12')
// (10, 22, 'sp12_v_b_11')
// (10, 23, 'sp12_v_b_8')
// (10, 24, 'sp12_v_b_7')
// (10, 25, 'sp12_v_b_4')
// (10, 26, 'sp12_v_b_3')
// (10, 27, 'sp12_h_l_23')
// (10, 27, 'sp12_v_b_0')
// (11, 15, 'sp4_h_r_21')
// (12, 15, 'sp4_h_r_32')
// (13, 15, 'sp4_h_r_45')
// (14, 15, 'sp4_h_l_45')
// (14, 15, 'sp4_h_r_8')
// (15, 15, 'local_g0_5')
// (15, 15, 'lutff_5/in_0')
// (15, 15, 'sp4_h_r_21')
// (16, 15, 'sp4_h_r_32')
// (16, 20, 'lutff_global/clk')
// (17, 15, 'sp4_h_r_45')
// (18, 15, 'sp4_h_l_45')
// (18, 23, 'lutff_global/clk')
// (24, 22, 'lutff_global/clk')
// (25, 15, 'ram/RCLK')
// (25, 17, 'ram/RCLK')
// (25, 19, 'ram/RCLK')
// (25, 21, 'ram/RCLK')
// (25, 23, 'ram/RCLK')
// (25, 25, 'ram/RCLK')
// (25, 27, 'ram/RCLK')
// (25, 29, 'ram/RCLK')

wire io_0_11_1;
assign io_0_11_1 = io_0_28_0;
// (0, 8, 'span4_vert_t_12')
// (0, 9, 'span4_vert_b_12')
// (0, 10, 'span4_vert_b_8')
// (0, 11, 'io_1/D_OUT_0')
// (0, 11, 'io_1/PAD')
// (0, 11, 'local_g1_4')
// (0, 11, 'span4_vert_b_4')
// (0, 12, 'span4_vert_b_0')
// (0, 12, 'span4_vert_t_12')
// (0, 13, 'span4_vert_b_12')
// (0, 14, 'span4_vert_b_8')
// (0, 15, 'span4_vert_b_4')
// (0, 16, 'span4_vert_b_0')
// (0, 16, 'span4_vert_t_12')
// (0, 17, 'span4_vert_b_12')
// (0, 18, 'span4_vert_b_8')
// (0, 19, 'span4_vert_b_4')
// (0, 20, 'span4_vert_b_0')
// (0, 20, 'span4_vert_t_12')
// (0, 21, 'span4_vert_b_12')
// (0, 22, 'span4_vert_b_8')
// (0, 23, 'span4_vert_b_4')
// (0, 24, 'span4_horz_25')
// (0, 24, 'span4_vert_b_0')
// (0, 24, 'span4_vert_t_12')
// (0, 25, 'span4_vert_b_12')
// (0, 26, 'span4_vert_b_8')
// (0, 27, 'span4_vert_b_4')
// (0, 28, 'io_0/D_IN_0')
// (0, 28, 'io_0/PAD')
// (0, 28, 'span4_vert_b_0')
// (1, 21, 'sp4_r_v_b_42')
// (1, 22, 'sp4_r_v_b_31')
// (1, 23, 'local_g3_2')
// (1, 23, 'lutff_0/in_1')
// (1, 23, 'sp4_r_v_b_18')
// (1, 24, 'sp4_h_r_36')
// (1, 24, 'sp4_r_v_b_7')
// (1, 27, 'neigh_op_tnl_0')
// (1, 27, 'neigh_op_tnl_4')
// (1, 28, 'neigh_op_lft_0')
// (1, 28, 'neigh_op_lft_4')
// (1, 29, 'neigh_op_bnl_0')
// (1, 29, 'neigh_op_bnl_4')
// (2, 20, 'sp4_v_t_42')
// (2, 21, 'sp4_v_b_42')
// (2, 22, 'sp4_v_b_31')
// (2, 23, 'sp4_v_b_18')
// (2, 24, 'sp4_h_l_36')
// (2, 24, 'sp4_v_b_7')

wire io_0_11_0;
// (0, 11, 'io_0/D_OUT_0')
// (0, 11, 'io_0/PAD')
// (0, 11, 'local_g1_5')
// (0, 11, 'span4_horz_5')
// (1, 11, 'sp4_h_r_16')
// (2, 11, 'sp4_h_r_29')
// (3, 11, 'sp4_h_r_40')
// (4, 11, 'sp4_h_l_40')
// (4, 11, 'sp4_h_r_5')
// (4, 20, 'sp4_h_r_5')
// (5, 11, 'sp4_h_r_16')
// (5, 20, 'sp4_h_r_16')
// (6, 11, 'sp4_h_r_29')
// (6, 20, 'local_g3_5')
// (6, 20, 'lutff_1/in_3')
// (6, 20, 'sp4_h_r_29')
// (7, 11, 'sp4_h_r_40')
// (7, 12, 'sp4_r_v_b_46')
// (7, 13, 'sp4_r_v_b_35')
// (7, 14, 'sp4_r_v_b_22')
// (7, 14, 'sp4_r_v_b_41')
// (7, 15, 'sp4_r_v_b_11')
// (7, 15, 'sp4_r_v_b_28')
// (7, 16, 'sp4_r_v_b_17')
// (7, 17, 'sp4_r_v_b_4')
// (7, 17, 'sp4_r_v_b_44')
// (7, 17, 'sp4_r_v_b_46')
// (7, 18, 'sp4_r_v_b_33')
// (7, 18, 'sp4_r_v_b_35')
// (7, 18, 'sp4_r_v_b_45')
// (7, 19, 'sp4_r_v_b_20')
// (7, 19, 'sp4_r_v_b_22')
// (7, 19, 'sp4_r_v_b_32')
// (7, 20, 'sp4_h_r_40')
// (7, 20, 'sp4_r_v_b_11')
// (7, 20, 'sp4_r_v_b_21')
// (7, 20, 'sp4_r_v_b_9')
// (7, 21, 'sp4_r_v_b_41')
// (7, 21, 'sp4_r_v_b_46')
// (7, 21, 'sp4_r_v_b_8')
// (7, 22, 'sp4_r_v_b_28')
// (7, 22, 'sp4_r_v_b_35')
// (7, 23, 'sp4_r_v_b_17')
// (7, 23, 'sp4_r_v_b_22')
// (7, 24, 'sp4_r_v_b_11')
// (7, 24, 'sp4_r_v_b_4')
// (7, 25, 'sp4_h_r_8')
// (7, 25, 'sp4_r_v_b_37')
// (7, 25, 'sp4_r_v_b_40')
// (7, 26, 'sp4_r_v_b_24')
// (7, 26, 'sp4_r_v_b_29')
// (7, 27, 'sp4_r_v_b_13')
// (7, 27, 'sp4_r_v_b_16')
// (7, 27, 'sp4_r_v_b_37')
// (7, 28, 'sp4_r_v_b_0')
// (7, 28, 'sp4_r_v_b_24')
// (7, 28, 'sp4_r_v_b_44')
// (7, 28, 'sp4_r_v_b_5')
// (7, 29, 'sp4_r_v_b_13')
// (7, 29, 'sp4_r_v_b_33')
// (7, 30, 'sp4_r_v_b_0')
// (7, 30, 'sp4_r_v_b_20')
// (7, 31, 'sp4_r_v_b_9')
// (8, 11, 'sp4_h_l_40')
// (8, 11, 'sp4_v_t_46')
// (8, 12, 'sp12_v_t_22')
// (8, 12, 'sp4_v_b_46')
// (8, 13, 'sp12_v_b_22')
// (8, 13, 'sp4_v_b_35')
// (8, 13, 'sp4_v_t_41')
// (8, 14, 'sp12_v_b_21')
// (8, 14, 'sp4_v_b_22')
// (8, 14, 'sp4_v_b_41')
// (8, 15, 'local_g2_4')
// (8, 15, 'ram/RE')
// (8, 15, 'sp12_v_b_18')
// (8, 15, 'sp4_v_b_11')
// (8, 15, 'sp4_v_b_28')
// (8, 16, 'local_g0_4')
// (8, 16, 'ram/WE')
// (8, 16, 'sp12_v_b_17')
// (8, 16, 'sp4_h_r_4')
// (8, 16, 'sp4_v_b_17')
// (8, 16, 'sp4_v_t_44')
// (8, 16, 'sp4_v_t_46')
// (8, 17, 'local_g1_5')
// (8, 17, 'ram/RE')
// (8, 17, 'sp12_v_b_14')
// (8, 17, 'sp4_h_r_11')
// (8, 17, 'sp4_h_r_5')
// (8, 17, 'sp4_v_b_4')
// (8, 17, 'sp4_v_b_44')
// (8, 17, 'sp4_v_b_46')
// (8, 17, 'sp4_v_t_45')
// (8, 18, 'local_g3_5')
// (8, 18, 'ram/WE')
// (8, 18, 'sp12_v_b_13')
// (8, 18, 'sp4_v_b_33')
// (8, 18, 'sp4_v_b_35')
// (8, 18, 'sp4_v_b_45')
// (8, 19, 'local_g0_4')
// (8, 19, 'ram/RE')
// (8, 19, 'sp12_v_b_10')
// (8, 19, 'sp4_v_b_20')
// (8, 19, 'sp4_v_b_22')
// (8, 19, 'sp4_v_b_32')
// (8, 20, 'local_g0_4')
// (8, 20, 'ram/WE')
// (8, 20, 'sp12_v_b_9')
// (8, 20, 'sp4_h_l_40')
// (8, 20, 'sp4_h_r_4')
// (8, 20, 'sp4_v_b_11')
// (8, 20, 'sp4_v_b_21')
// (8, 20, 'sp4_v_b_9')
// (8, 20, 'sp4_v_t_41')
// (8, 20, 'sp4_v_t_46')
// (8, 21, 'local_g1_5')
// (8, 21, 'ram/RE')
// (8, 21, 'sp12_v_b_6')
// (8, 21, 'sp4_h_r_5')
// (8, 21, 'sp4_h_r_8')
// (8, 21, 'sp4_v_b_41')
// (8, 21, 'sp4_v_b_46')
// (8, 21, 'sp4_v_b_8')
// (8, 22, 'local_g2_4')
// (8, 22, 'ram/WE')
// (8, 22, 'sp12_v_b_5')
// (8, 22, 'sp4_v_b_28')
// (8, 22, 'sp4_v_b_35')
// (8, 23, 'local_g0_4')
// (8, 23, 'ram/RE')
// (8, 23, 'sp12_v_b_2')
// (8, 23, 'sp4_h_r_4')
// (8, 23, 'sp4_v_b_17')
// (8, 23, 'sp4_v_b_22')
// (8, 24, 'local_g0_4')
// (8, 24, 'ram/WE')
// (8, 24, 'sp12_h_r_1')
// (8, 24, 'sp12_v_b_1')
// (8, 24, 'sp4_h_r_11')
// (8, 24, 'sp4_v_b_11')
// (8, 24, 'sp4_v_b_4')
// (8, 24, 'sp4_v_t_37')
// (8, 24, 'sp4_v_t_40')
// (8, 25, 'local_g1_5')
// (8, 25, 'ram/RE')
// (8, 25, 'sp4_h_r_21')
// (8, 25, 'sp4_v_b_37')
// (8, 25, 'sp4_v_b_40')
// (8, 26, 'local_g3_5')
// (8, 26, 'ram/WE')
// (8, 26, 'sp4_h_r_0')
// (8, 26, 'sp4_v_b_24')
// (8, 26, 'sp4_v_b_29')
// (8, 26, 'sp4_v_t_37')
// (8, 27, 'local_g1_5')
// (8, 27, 'ram/RE')
// (8, 27, 'sp4_h_r_3')
// (8, 27, 'sp4_v_b_13')
// (8, 27, 'sp4_v_b_16')
// (8, 27, 'sp4_v_b_37')
// (8, 27, 'sp4_v_t_44')
// (8, 28, 'local_g1_5')
// (8, 28, 'ram/WE')
// (8, 28, 'sp4_v_b_0')
// (8, 28, 'sp4_v_b_24')
// (8, 28, 'sp4_v_b_44')
// (8, 28, 'sp4_v_b_5')
// (8, 29, 'local_g1_5')
// (8, 29, 'ram/RE')
// (8, 29, 'sp4_v_b_13')
// (8, 29, 'sp4_v_b_33')
// (8, 30, 'local_g0_4')
// (8, 30, 'ram/WE')
// (8, 30, 'sp4_v_b_0')
// (8, 30, 'sp4_v_b_20')
// (8, 31, 'sp4_v_b_9')
// (9, 16, 'sp4_h_r_17')
// (9, 17, 'sp4_h_r_16')
// (9, 17, 'sp4_h_r_22')
// (9, 20, 'sp4_h_r_17')
// (9, 21, 'sp4_h_r_16')
// (9, 21, 'sp4_h_r_21')
// (9, 23, 'sp4_h_r_17')
// (9, 24, 'sp12_h_r_2')
// (9, 24, 'sp4_h_r_22')
// (9, 25, 'sp4_h_r_32')
// (9, 26, 'sp4_h_r_13')
// (9, 27, 'sp4_h_r_14')
// (10, 16, 'sp4_h_r_28')
// (10, 17, 'sp4_h_r_29')
// (10, 17, 'sp4_h_r_35')
// (10, 20, 'sp4_h_r_28')
// (10, 21, 'sp4_h_r_29')
// (10, 21, 'sp4_h_r_32')
// (10, 22, 'sp4_r_v_b_38')
// (10, 23, 'neigh_op_tnr_7')
// (10, 23, 'sp4_h_r_28')
// (10, 23, 'sp4_r_v_b_27')
// (10, 24, 'neigh_op_rgt_7')
// (10, 24, 'sp12_h_r_5')
// (10, 24, 'sp4_h_r_3')
// (10, 24, 'sp4_h_r_35')
// (10, 24, 'sp4_r_v_b_14')
// (10, 25, 'neigh_op_bnr_7')
// (10, 25, 'sp4_h_r_45')
// (10, 25, 'sp4_r_v_b_3')
// (10, 26, 'sp4_h_r_24')
// (10, 27, 'sp4_h_r_27')
// (11, 16, 'sp4_h_r_41')
// (11, 17, 'sp4_h_r_40')
// (11, 17, 'sp4_h_r_46')
// (11, 18, 'sp4_r_v_b_40')
// (11, 19, 'sp4_r_v_b_29')
// (11, 20, 'sp4_h_r_41')
// (11, 20, 'sp4_r_v_b_16')
// (11, 21, 'sp4_h_r_40')
// (11, 21, 'sp4_h_r_45')
// (11, 21, 'sp4_r_v_b_5')
// (11, 21, 'sp4_v_t_38')
// (11, 22, 'sp4_r_v_b_39')
// (11, 22, 'sp4_v_b_38')
// (11, 23, 'neigh_op_top_7')
// (11, 23, 'sp4_h_r_41')
// (11, 23, 'sp4_r_v_b_26')
// (11, 23, 'sp4_r_v_b_42')
// (11, 23, 'sp4_v_b_27')
// (11, 24, 'lutff_7/out')
// (11, 24, 'sp12_h_r_6')
// (11, 24, 'sp4_h_r_14')
// (11, 24, 'sp4_h_r_46')
// (11, 24, 'sp4_r_v_b_15')
// (11, 24, 'sp4_r_v_b_31')
// (11, 24, 'sp4_r_v_b_47')
// (11, 24, 'sp4_v_b_14')
// (11, 25, 'neigh_op_bot_7')
// (11, 25, 'sp4_h_l_45')
// (11, 25, 'sp4_r_v_b_18')
// (11, 25, 'sp4_r_v_b_2')
// (11, 25, 'sp4_r_v_b_34')
// (11, 25, 'sp4_v_b_3')
// (11, 26, 'sp4_h_r_37')
// (11, 26, 'sp4_r_v_b_23')
// (11, 26, 'sp4_r_v_b_7')
// (11, 27, 'sp4_h_r_38')
// (11, 27, 'sp4_r_v_b_10')
// (12, 16, 'sp4_h_l_41')
// (12, 17, 'sp4_h_l_40')
// (12, 17, 'sp4_h_l_46')
// (12, 17, 'sp4_v_t_40')
// (12, 18, 'sp4_v_b_40')
// (12, 19, 'sp4_v_b_29')
// (12, 20, 'sp4_h_l_41')
// (12, 20, 'sp4_v_b_16')
// (12, 21, 'sp4_h_l_40')
// (12, 21, 'sp4_h_l_45')
// (12, 21, 'sp4_h_r_2')
// (12, 21, 'sp4_h_r_7')
// (12, 21, 'sp4_v_b_5')
// (12, 21, 'sp4_v_t_39')
// (12, 22, 'sp4_v_b_39')
// (12, 22, 'sp4_v_t_42')
// (12, 23, 'neigh_op_tnl_7')
// (12, 23, 'sp4_h_l_41')
// (12, 23, 'sp4_v_b_26')
// (12, 23, 'sp4_v_b_42')
// (12, 23, 'sp4_v_t_47')
// (12, 24, 'neigh_op_lft_7')
// (12, 24, 'sp12_h_r_9')
// (12, 24, 'sp4_h_l_46')
// (12, 24, 'sp4_h_r_27')
// (12, 24, 'sp4_v_b_15')
// (12, 24, 'sp4_v_b_31')
// (12, 24, 'sp4_v_b_47')
// (12, 25, 'neigh_op_bnl_7')
// (12, 25, 'sp4_h_r_2')
// (12, 25, 'sp4_v_b_18')
// (12, 25, 'sp4_v_b_2')
// (12, 25, 'sp4_v_b_34')
// (12, 26, 'sp4_h_l_37')
// (12, 26, 'sp4_h_r_1')
// (12, 26, 'sp4_v_b_23')
// (12, 26, 'sp4_v_b_7')
// (12, 27, 'sp4_h_l_38')
// (12, 27, 'sp4_v_b_10')
// (13, 13, 'sp4_r_v_b_38')
// (13, 14, 'sp4_r_v_b_27')
// (13, 15, 'sp4_r_v_b_14')
// (13, 16, 'sp4_r_v_b_3')
// (13, 17, 'sp4_r_v_b_38')
// (13, 18, 'sp4_r_v_b_27')
// (13, 19, 'sp4_r_v_b_14')
// (13, 20, 'sp4_r_v_b_3')
// (13, 21, 'sp4_h_r_15')
// (13, 21, 'sp4_h_r_18')
// (13, 21, 'sp4_r_v_b_38')
// (13, 22, 'sp4_r_v_b_27')
// (13, 23, 'sp4_r_v_b_14')
// (13, 24, 'sp12_h_r_10')
// (13, 24, 'sp4_h_r_38')
// (13, 24, 'sp4_r_v_b_3')
// (13, 25, 'sp4_h_r_15')
// (13, 26, 'sp4_h_r_12')
// (14, 12, 'sp4_h_r_3')
// (14, 12, 'sp4_v_t_38')
// (14, 13, 'sp4_v_b_38')
// (14, 14, 'sp4_v_b_27')
// (14, 15, 'sp4_v_b_14')
// (14, 16, 'sp4_h_r_8')
// (14, 16, 'sp4_v_b_3')
// (14, 16, 'sp4_v_t_38')
// (14, 17, 'sp4_v_b_38')
// (14, 18, 'sp4_v_b_27')
// (14, 19, 'sp4_v_b_14')
// (14, 20, 'sp4_h_r_8')
// (14, 20, 'sp4_v_b_3')
// (14, 20, 'sp4_v_t_38')
// (14, 21, 'sp4_h_r_26')
// (14, 21, 'sp4_h_r_31')
// (14, 21, 'sp4_v_b_38')
// (14, 22, 'sp4_v_b_27')
// (14, 23, 'sp4_v_b_14')
// (14, 24, 'sp12_h_r_13')
// (14, 24, 'sp4_h_l_38')
// (14, 24, 'sp4_h_r_6')
// (14, 24, 'sp4_v_b_3')
// (14, 25, 'sp4_h_r_26')
// (14, 26, 'sp4_h_r_25')
// (15, 10, 'sp4_r_v_b_37')
// (15, 11, 'sp4_r_v_b_24')
// (15, 12, 'sp4_h_r_14')
// (15, 12, 'sp4_r_v_b_13')
// (15, 13, 'sp4_r_v_b_0')
// (15, 14, 'sp4_r_v_b_41')
// (15, 15, 'sp4_r_v_b_28')
// (15, 16, 'sp4_h_r_21')
// (15, 16, 'sp4_r_v_b_17')
// (15, 17, 'sp4_r_v_b_4')
// (15, 18, 'sp4_r_v_b_36')
// (15, 19, 'sp4_r_v_b_25')
// (15, 20, 'sp4_h_r_21')
// (15, 20, 'sp4_r_v_b_12')
// (15, 21, 'sp4_h_r_39')
// (15, 21, 'sp4_h_r_42')
// (15, 21, 'sp4_r_v_b_1')
// (15, 24, 'sp12_h_r_14')
// (15, 24, 'sp4_h_r_19')
// (15, 25, 'sp4_h_r_39')
// (15, 26, 'sp4_h_r_36')
// (16, 9, 'sp4_v_t_37')
// (16, 10, 'sp4_v_b_37')
// (16, 11, 'local_g2_0')
// (16, 11, 'local_g3_0')
// (16, 11, 'lutff_1/in_1')
// (16, 11, 'lutff_2/in_2')
// (16, 11, 'lutff_3/in_2')
// (16, 11, 'lutff_4/in_2')
// (16, 11, 'lutff_5/in_1')
// (16, 11, 'lutff_6/in_2')
// (16, 11, 'lutff_7/in_2')
// (16, 11, 'sp4_v_b_24')
// (16, 12, 'local_g0_5')
// (16, 12, 'local_g1_5')
// (16, 12, 'lutff_0/in_1')
// (16, 12, 'lutff_1/in_2')
// (16, 12, 'lutff_2/in_2')
// (16, 12, 'lutff_3/in_2')
// (16, 12, 'lutff_4/in_1')
// (16, 12, 'lutff_5/in_2')
// (16, 12, 'lutff_6/in_2')
// (16, 12, 'lutff_7/in_0')
// (16, 12, 'sp4_h_r_27')
// (16, 12, 'sp4_v_b_13')
// (16, 13, 'sp4_v_b_0')
// (16, 13, 'sp4_v_t_41')
// (16, 14, 'local_g2_1')
// (16, 14, 'lutff_3/in_2')
// (16, 14, 'sp4_v_b_41')
// (16, 15, 'sp4_v_b_28')
// (16, 16, 'sp4_h_r_32')
// (16, 16, 'sp4_v_b_17')
// (16, 17, 'sp4_v_b_4')
// (16, 17, 'sp4_v_t_36')
// (16, 18, 'sp4_v_b_36')
// (16, 19, 'sp4_v_b_25')
// (16, 20, 'sp4_h_r_32')
// (16, 20, 'sp4_v_b_12')
// (16, 21, 'sp4_h_l_39')
// (16, 21, 'sp4_h_l_42')
// (16, 21, 'sp4_h_r_3')
// (16, 21, 'sp4_v_b_1')
// (16, 24, 'sp12_h_r_17')
// (16, 24, 'sp4_h_r_30')
// (16, 25, 'sp4_h_l_39')
// (16, 25, 'sp4_h_r_10')
// (16, 25, 'sp4_h_r_5')
// (16, 26, 'sp4_h_l_36')
// (16, 26, 'sp4_h_r_9')
// (17, 9, 'sp4_r_v_b_38')
// (17, 10, 'sp4_r_v_b_27')
// (17, 11, 'local_g2_6')
// (17, 11, 'lutff_7/in_1')
// (17, 11, 'sp4_r_v_b_14')
// (17, 12, 'sp4_h_r_38')
// (17, 12, 'sp4_r_v_b_3')
// (17, 16, 'sp4_h_r_45')
// (17, 20, 'sp4_h_r_45')
// (17, 21, 'sp4_h_r_14')
// (17, 24, 'sp12_h_r_18')
// (17, 24, 'sp4_h_r_43')
// (17, 25, 'sp4_h_r_16')
// (17, 25, 'sp4_h_r_23')
// (17, 26, 'sp4_h_r_20')
// (18, 8, 'sp4_v_t_38')
// (18, 9, 'sp4_v_b_38')
// (18, 10, 'sp4_v_b_27')
// (18, 11, 'sp4_v_b_14')
// (18, 12, 'sp4_h_l_38')
// (18, 12, 'sp4_v_b_3')
// (18, 16, 'sp4_h_l_45')
// (18, 16, 'sp4_h_r_4')
// (18, 20, 'sp4_h_l_45')
// (18, 20, 'sp4_h_r_8')
// (18, 21, 'sp4_h_r_27')
// (18, 24, 'sp12_h_r_21')
// (18, 24, 'sp4_h_l_43')
// (18, 24, 'sp4_h_r_2')
// (18, 25, 'sp4_h_r_29')
// (18, 25, 'sp4_h_r_34')
// (18, 26, 'sp4_h_r_33')
// (19, 12, 'sp4_r_v_b_46')
// (19, 13, 'sp4_r_v_b_35')
// (19, 14, 'sp4_r_v_b_22')
// (19, 15, 'sp4_r_v_b_11')
// (19, 16, 'sp4_h_r_17')
// (19, 18, 'sp4_r_v_b_44')
// (19, 19, 'sp4_r_v_b_33')
// (19, 20, 'sp4_h_r_21')
// (19, 20, 'sp4_r_v_b_20')
// (19, 21, 'sp4_h_r_38')
// (19, 21, 'sp4_r_v_b_9')
// (19, 24, 'sp12_h_r_22')
// (19, 24, 'sp4_h_r_15')
// (19, 25, 'sp4_h_r_40')
// (19, 25, 'sp4_h_r_47')
// (19, 26, 'sp4_h_r_44')
// (20, 11, 'sp4_v_t_46')
// (20, 12, 'sp12_v_t_22')
// (20, 12, 'sp4_v_b_46')
// (20, 13, 'sp12_v_b_22')
// (20, 13, 'sp4_v_b_35')
// (20, 14, 'sp12_v_b_21')
// (20, 14, 'sp4_v_b_22')
// (20, 15, 'sp12_v_b_18')
// (20, 15, 'sp4_h_r_5')
// (20, 15, 'sp4_v_b_11')
// (20, 16, 'sp12_v_b_17')
// (20, 16, 'sp4_h_r_28')
// (20, 17, 'sp12_v_b_14')
// (20, 17, 'sp4_h_r_9')
// (20, 17, 'sp4_v_t_44')
// (20, 18, 'sp12_v_b_13')
// (20, 18, 'sp4_v_b_44')
// (20, 19, 'sp12_v_b_10')
// (20, 19, 'sp4_v_b_33')
// (20, 20, 'sp12_v_b_9')
// (20, 20, 'sp4_h_r_32')
// (20, 20, 'sp4_v_b_20')
// (20, 21, 'sp12_v_b_6')
// (20, 21, 'sp4_h_l_38')
// (20, 21, 'sp4_h_r_6')
// (20, 21, 'sp4_v_b_9')
// (20, 22, 'sp12_v_b_5')
// (20, 23, 'sp12_v_b_2')
// (20, 24, 'sp12_h_l_22')
// (20, 24, 'sp12_v_b_1')
// (20, 24, 'sp4_h_r_26')
// (20, 25, 'sp4_h_l_40')
// (20, 25, 'sp4_h_l_47')
// (20, 25, 'sp4_h_r_5')
// (20, 25, 'sp4_h_r_6')
// (20, 26, 'sp4_h_l_44')
// (20, 26, 'sp4_h_r_0')
// (21, 15, 'sp4_h_r_16')
// (21, 16, 'sp4_h_r_41')
// (21, 17, 'sp4_h_r_20')
// (21, 20, 'local_g2_5')
// (21, 20, 'lutff_5/in_2')
// (21, 20, 'sp4_h_r_45')
// (21, 21, 'sp4_h_r_19')
// (21, 24, 'sp4_h_r_39')
// (21, 25, 'sp4_h_r_16')
// (21, 25, 'sp4_h_r_19')
// (21, 26, 'sp4_h_r_13')
// (22, 15, 'sp4_h_r_29')
// (22, 16, 'sp4_h_l_41')
// (22, 16, 'sp4_h_r_0')
// (22, 17, 'sp4_h_r_33')
// (22, 20, 'sp4_h_l_45')
// (22, 20, 'sp4_h_r_11')
// (22, 20, 'sp4_h_r_8')
// (22, 21, 'sp4_h_r_30')
// (22, 24, 'sp4_h_l_39')
// (22, 24, 'sp4_h_r_2')
// (22, 24, 'sp4_h_r_5')
// (22, 25, 'sp4_h_r_29')
// (22, 25, 'sp4_h_r_30')
// (22, 26, 'sp4_h_r_24')
// (23, 15, 'sp4_h_r_40')
// (23, 16, 'sp4_h_r_13')
// (23, 17, 'sp4_h_r_44')
// (23, 18, 'sp4_r_v_b_43')
// (23, 19, 'sp4_r_v_b_30')
// (23, 20, 'sp4_h_r_21')
// (23, 20, 'sp4_h_r_22')
// (23, 20, 'sp4_r_v_b_19')
// (23, 21, 'sp4_h_r_43')
// (23, 21, 'sp4_r_v_b_6')
// (23, 24, 'sp4_h_r_15')
// (23, 24, 'sp4_h_r_16')
// (23, 25, 'sp4_h_r_40')
// (23, 25, 'sp4_h_r_43')
// (23, 26, 'sp4_h_r_37')
// (23, 26, 'sp4_r_v_b_43')
// (23, 27, 'sp4_r_v_b_30')
// (23, 27, 'sp4_r_v_b_37')
// (23, 28, 'sp4_r_v_b_19')
// (23, 28, 'sp4_r_v_b_24')
// (23, 29, 'sp4_r_v_b_13')
// (23, 29, 'sp4_r_v_b_6')
// (23, 30, 'sp4_r_v_b_0')
// (24, 15, 'sp4_h_l_40')
// (24, 15, 'sp4_h_r_1')
// (24, 16, 'sp4_h_r_24')
// (24, 17, 'sp4_h_l_44')
// (24, 17, 'sp4_h_r_0')
// (24, 17, 'sp4_v_t_43')
// (24, 18, 'sp4_v_b_43')
// (24, 19, 'sp4_v_b_30')
// (24, 20, 'sp4_h_r_32')
// (24, 20, 'sp4_h_r_35')
// (24, 20, 'sp4_v_b_19')
// (24, 21, 'sp4_h_l_43')
// (24, 21, 'sp4_h_r_0')
// (24, 21, 'sp4_v_b_6')
// (24, 24, 'sp4_h_r_26')
// (24, 24, 'sp4_h_r_29')
// (24, 25, 'sp4_h_l_40')
// (24, 25, 'sp4_h_l_43')
// (24, 25, 'sp4_h_r_8')
// (24, 25, 'sp4_v_t_43')
// (24, 26, 'sp4_h_l_37')
// (24, 26, 'sp4_v_b_43')
// (24, 26, 'sp4_v_t_37')
// (24, 27, 'sp4_v_b_30')
// (24, 27, 'sp4_v_b_37')
// (24, 28, 'sp4_v_b_19')
// (24, 28, 'sp4_v_b_24')
// (24, 29, 'sp4_h_r_0')
// (24, 29, 'sp4_v_b_13')
// (24, 29, 'sp4_v_b_6')
// (24, 30, 'sp4_h_r_0')
// (24, 30, 'sp4_v_b_0')
// (25, 15, 'local_g0_4')
// (25, 15, 'ram/RE')
// (25, 15, 'sp4_h_r_12')
// (25, 16, 'local_g3_5')
// (25, 16, 'ram/WE')
// (25, 16, 'sp4_h_r_37')
// (25, 17, 'local_g1_5')
// (25, 17, 'ram/RE')
// (25, 17, 'sp4_h_r_13')
// (25, 17, 'sp4_r_v_b_40')
// (25, 17, 'sp4_r_v_b_45')
// (25, 18, 'local_g1_5')
// (25, 18, 'ram/WE')
// (25, 18, 'sp4_r_v_b_29')
// (25, 18, 'sp4_r_v_b_32')
// (25, 19, 'local_g3_5')
// (25, 19, 'ram/RE')
// (25, 19, 'sp4_r_v_b_16')
// (25, 19, 'sp4_r_v_b_21')
// (25, 20, 'local_g3_5')
// (25, 20, 'ram/WE')
// (25, 20, 'sp4_h_r_45')
// (25, 20, 'sp4_h_r_46')
// (25, 20, 'sp4_r_v_b_5')
// (25, 20, 'sp4_r_v_b_8')
// (25, 21, 'local_g1_5')
// (25, 21, 'ram/RE')
// (25, 21, 'sp4_h_r_13')
// (25, 21, 'sp4_r_v_b_40')
// (25, 21, 'sp4_r_v_b_45')
// (25, 22, 'local_g1_5')
// (25, 22, 'ram/WE')
// (25, 22, 'sp4_r_v_b_29')
// (25, 22, 'sp4_r_v_b_32')
// (25, 23, 'local_g3_5')
// (25, 23, 'ram/RE')
// (25, 23, 'sp4_r_v_b_16')
// (25, 23, 'sp4_r_v_b_21')
// (25, 24, 'local_g1_5')
// (25, 24, 'ram/WE')
// (25, 24, 'sp4_h_r_39')
// (25, 24, 'sp4_h_r_40')
// (25, 24, 'sp4_r_v_b_5')
// (25, 24, 'sp4_r_v_b_8')
// (25, 25, 'local_g1_5')
// (25, 25, 'ram/RE')
// (25, 25, 'sp4_h_r_21')
// (25, 25, 'sp4_r_v_b_40')
// (25, 25, 'sp4_r_v_b_45')
// (25, 26, 'local_g1_5')
// (25, 26, 'ram/WE')
// (25, 26, 'sp4_r_v_b_29')
// (25, 26, 'sp4_r_v_b_32')
// (25, 27, 'local_g3_5')
// (25, 27, 'ram/RE')
// (25, 27, 'sp4_r_v_b_16')
// (25, 27, 'sp4_r_v_b_21')
// (25, 28, 'local_g1_5')
// (25, 28, 'ram/WE')
// (25, 28, 'sp4_r_v_b_5')
// (25, 28, 'sp4_r_v_b_8')
// (25, 29, 'local_g1_5')
// (25, 29, 'ram/RE')
// (25, 29, 'sp4_h_r_13')
// (25, 30, 'local_g1_5')
// (25, 30, 'ram/WE')
// (25, 30, 'sp4_h_r_13')
// (26, 15, 'sp4_h_r_25')
// (26, 16, 'sp4_h_l_37')
// (26, 16, 'sp4_v_t_40')
// (26, 16, 'sp4_v_t_45')
// (26, 17, 'sp4_h_r_24')
// (26, 17, 'sp4_v_b_40')
// (26, 17, 'sp4_v_b_45')
// (26, 18, 'sp4_v_b_29')
// (26, 18, 'sp4_v_b_32')
// (26, 19, 'sp4_v_b_16')
// (26, 19, 'sp4_v_b_21')
// (26, 20, 'sp4_h_l_45')
// (26, 20, 'sp4_h_l_46')
// (26, 20, 'sp4_v_b_5')
// (26, 20, 'sp4_v_b_8')
// (26, 20, 'sp4_v_t_40')
// (26, 20, 'sp4_v_t_45')
// (26, 21, 'sp4_h_r_24')
// (26, 21, 'sp4_v_b_40')
// (26, 21, 'sp4_v_b_45')
// (26, 22, 'sp4_v_b_29')
// (26, 22, 'sp4_v_b_32')
// (26, 23, 'sp4_v_b_16')
// (26, 23, 'sp4_v_b_21')
// (26, 24, 'sp4_h_l_39')
// (26, 24, 'sp4_h_l_40')
// (26, 24, 'sp4_h_r_8')
// (26, 24, 'sp4_v_b_5')
// (26, 24, 'sp4_v_b_8')
// (26, 24, 'sp4_v_t_40')
// (26, 24, 'sp4_v_t_45')
// (26, 25, 'sp4_h_r_32')
// (26, 25, 'sp4_v_b_40')
// (26, 25, 'sp4_v_b_45')
// (26, 26, 'sp4_v_b_29')
// (26, 26, 'sp4_v_b_32')
// (26, 27, 'sp4_v_b_16')
// (26, 27, 'sp4_v_b_21')
// (26, 28, 'sp4_v_b_5')
// (26, 28, 'sp4_v_b_8')
// (26, 29, 'sp4_h_r_24')
// (26, 30, 'sp4_h_r_24')
// (27, 15, 'sp4_h_r_36')
// (27, 17, 'sp4_h_r_37')
// (27, 21, 'sp4_h_r_37')
// (27, 24, 'sp4_h_r_21')
// (27, 25, 'sp4_h_r_45')
// (27, 29, 'sp4_h_r_37')
// (27, 30, 'sp4_h_r_37')
// (28, 15, 'sp4_h_l_36')
// (28, 17, 'sp4_h_l_37')
// (28, 21, 'sp4_h_l_37')
// (28, 24, 'sp4_h_r_32')
// (28, 25, 'sp4_h_l_45')
// (28, 29, 'sp4_h_l_37')
// (28, 30, 'sp4_h_l_37')
// (29, 24, 'sp4_h_r_45')
// (30, 24, 'sp4_h_l_45')

reg io_0_18_1 = 0;
// (0, 15, 'span4_vert_t_12')
// (0, 16, 'span4_vert_b_12')
// (0, 17, 'span4_vert_b_8')
// (0, 18, 'io_1/D_OUT_0')
// (0, 18, 'io_1/PAD')
// (0, 18, 'local_g1_4')
// (0, 18, 'span4_vert_b_4')
// (0, 19, 'span4_horz_25')
// (0, 19, 'span4_vert_b_0')
// (1, 19, 'sp4_h_r_36')
// (2, 19, 'sp4_h_l_36')
// (2, 19, 'sp4_h_r_5')
// (3, 19, 'sp4_h_r_16')
// (4, 19, 'sp4_h_r_29')
// (5, 19, 'sp4_h_r_40')
// (6, 18, 'neigh_op_tnr_0')
// (6, 19, 'neigh_op_rgt_0')
// (6, 19, 'sp4_h_l_40')
// (6, 19, 'sp4_h_r_5')
// (6, 20, 'neigh_op_bnr_0')
// (7, 18, 'neigh_op_top_0')
// (7, 19, 'lutff_0/out')
// (7, 19, 'sp4_h_r_16')
// (7, 20, 'neigh_op_bot_0')
// (8, 18, 'neigh_op_tnl_0')
// (8, 19, 'neigh_op_lft_0')
// (8, 19, 'sp4_h_r_29')
// (8, 20, 'neigh_op_bnl_0')
// (9, 19, 'sp4_h_r_40')
// (10, 19, 'sp4_h_l_40')

reg io_0_17_1 = 0;
// (0, 15, 'span4_vert_t_13')
// (0, 16, 'span4_vert_b_13')
// (0, 17, 'io_1/D_OUT_0')
// (0, 17, 'io_1/PAD')
// (0, 17, 'local_g0_1')
// (0, 17, 'span4_vert_b_9')
// (0, 18, 'span4_vert_b_5')
// (0, 19, 'span4_horz_31')
// (0, 19, 'span4_vert_b_1')
// (1, 19, 'sp4_h_r_42')
// (2, 19, 'sp4_h_l_42')
// (2, 19, 'sp4_h_r_7')
// (3, 19, 'sp4_h_r_18')
// (4, 19, 'sp4_h_r_31')
// (5, 19, 'sp4_h_r_42')
// (6, 18, 'neigh_op_tnr_3')
// (6, 19, 'neigh_op_rgt_3')
// (6, 19, 'sp4_h_l_42')
// (6, 19, 'sp4_h_r_11')
// (6, 20, 'neigh_op_bnr_3')
// (7, 18, 'neigh_op_top_3')
// (7, 19, 'lutff_3/out')
// (7, 19, 'sp4_h_r_22')
// (7, 20, 'neigh_op_bot_3')
// (8, 18, 'neigh_op_tnl_3')
// (8, 19, 'neigh_op_lft_3')
// (8, 19, 'sp4_h_r_35')
// (8, 20, 'neigh_op_bnl_3')
// (9, 19, 'sp4_h_r_46')
// (10, 19, 'sp4_h_l_46')

reg io_0_17_0 = 0;
// (0, 17, 'io_0/D_OUT_0')
// (0, 17, 'io_0/PAD')
// (0, 17, 'local_g0_2')
// (0, 17, 'span4_horz_18')
// (1, 17, 'sp4_h_r_31')
// (2, 17, 'sp4_h_r_42')
// (3, 17, 'sp4_h_l_42')
// (3, 17, 'sp4_h_r_4')
// (4, 17, 'sp4_h_r_17')
// (5, 17, 'sp4_h_r_28')
// (6, 17, 'sp4_h_r_41')
// (6, 18, 'sp4_r_v_b_47')
// (6, 19, 'sp4_r_v_b_34')
// (6, 20, 'neigh_op_tnr_5')
// (6, 20, 'sp4_r_v_b_23')
// (6, 21, 'neigh_op_rgt_5')
// (6, 21, 'sp4_r_v_b_10')
// (6, 22, 'neigh_op_bnr_5')
// (7, 17, 'sp4_h_l_41')
// (7, 17, 'sp4_v_t_47')
// (7, 18, 'sp4_v_b_47')
// (7, 19, 'sp4_v_b_34')
// (7, 20, 'neigh_op_top_5')
// (7, 20, 'sp4_v_b_23')
// (7, 21, 'lutff_5/out')
// (7, 21, 'sp4_v_b_10')
// (7, 22, 'neigh_op_bot_5')
// (8, 20, 'neigh_op_tnl_5')
// (8, 21, 'neigh_op_lft_5')
// (8, 22, 'neigh_op_bnl_5')

wire io_33_29_1;
// (0, 17, 'span12_horz_4')
// (1, 17, 'sp12_h_r_7')
// (2, 17, 'sp12_h_r_8')
// (3, 17, 'sp12_h_r_11')
// (4, 17, 'sp12_h_r_12')
// (5, 17, 'sp12_h_r_15')
// (6, 15, 'sp4_h_r_4')
// (6, 17, 'sp12_h_r_16')
// (6, 19, 'sp4_h_r_3')
// (6, 21, 'sp4_h_r_4')
// (7, 15, 'sp4_h_r_17')
// (7, 17, 'sp12_h_r_19')
// (7, 19, 'sp4_h_r_14')
// (7, 21, 'sp4_h_r_17')
// (7, 29, 'sp4_h_r_6')
// (8, 15, 'local_g3_4')
// (8, 15, 'ram/RADDR_8')
// (8, 15, 'sp4_h_r_28')
// (8, 17, 'local_g1_4')
// (8, 17, 'ram/RADDR_8')
// (8, 17, 'sp12_h_r_20')
// (8, 19, 'local_g2_3')
// (8, 19, 'ram/RADDR_8')
// (8, 19, 'sp4_h_r_27')
// (8, 21, 'local_g3_4')
// (8, 21, 'ram/RADDR_8')
// (8, 21, 'sp4_h_r_28')
// (8, 22, 'sp4_r_v_b_39')
// (8, 23, 'local_g1_2')
// (8, 23, 'ram/RADDR_8')
// (8, 23, 'sp4_r_v_b_26')
// (8, 24, 'sp4_r_v_b_15')
// (8, 25, 'local_g1_2')
// (8, 25, 'ram/RADDR_8')
// (8, 25, 'sp4_r_v_b_2')
// (8, 26, 'sp4_r_v_b_36')
// (8, 26, 'sp4_r_v_b_43')
// (8, 27, 'local_g0_1')
// (8, 27, 'ram/RADDR_8')
// (8, 27, 'sp4_r_v_b_25')
// (8, 27, 'sp4_r_v_b_30')
// (8, 28, 'sp4_r_v_b_12')
// (8, 28, 'sp4_r_v_b_19')
// (8, 29, 'local_g0_3')
// (8, 29, 'ram/RADDR_8')
// (8, 29, 'sp4_h_r_19')
// (8, 29, 'sp4_r_v_b_1')
// (8, 29, 'sp4_r_v_b_6')
// (9, 15, 'sp4_h_r_41')
// (9, 16, 'sp4_r_v_b_47')
// (9, 17, 'sp12_h_r_23')
// (9, 17, 'sp4_r_v_b_34')
// (9, 18, 'sp4_r_v_b_23')
// (9, 19, 'sp4_h_r_38')
// (9, 19, 'sp4_r_v_b_10')
// (9, 21, 'sp4_h_r_41')
// (9, 21, 'sp4_v_t_39')
// (9, 22, 'sp4_r_v_b_41')
// (9, 22, 'sp4_v_b_39')
// (9, 23, 'sp4_r_v_b_28')
// (9, 23, 'sp4_v_b_26')
// (9, 24, 'sp4_r_v_b_17')
// (9, 24, 'sp4_v_b_15')
// (9, 25, 'sp4_r_v_b_4')
// (9, 25, 'sp4_v_b_2')
// (9, 25, 'sp4_v_t_36')
// (9, 25, 'sp4_v_t_43')
// (9, 26, 'sp4_v_b_36')
// (9, 26, 'sp4_v_b_43')
// (9, 27, 'sp4_v_b_25')
// (9, 27, 'sp4_v_b_30')
// (9, 28, 'sp4_v_b_12')
// (9, 28, 'sp4_v_b_19')
// (9, 29, 'sp4_h_r_1')
// (9, 29, 'sp4_h_r_30')
// (9, 29, 'sp4_v_b_1')
// (9, 29, 'sp4_v_b_6')
// (10, 15, 'sp4_h_l_41')
// (10, 15, 'sp4_v_t_47')
// (10, 16, 'sp4_v_b_47')
// (10, 17, 'sp12_h_l_23')
// (10, 17, 'sp12_v_t_23')
// (10, 17, 'sp4_v_b_34')
// (10, 18, 'sp12_v_b_23')
// (10, 18, 'sp4_v_b_23')
// (10, 19, 'sp12_v_b_20')
// (10, 19, 'sp4_h_l_38')
// (10, 19, 'sp4_v_b_10')
// (10, 20, 'sp12_v_b_19')
// (10, 21, 'sp12_v_b_16')
// (10, 21, 'sp4_h_l_41')
// (10, 21, 'sp4_v_t_41')
// (10, 22, 'sp12_v_b_15')
// (10, 22, 'sp4_v_b_41')
// (10, 23, 'sp12_v_b_12')
// (10, 23, 'sp4_v_b_28')
// (10, 24, 'sp12_v_b_11')
// (10, 24, 'sp4_v_b_17')
// (10, 25, 'sp12_v_b_8')
// (10, 25, 'sp4_v_b_4')
// (10, 26, 'sp12_v_b_7')
// (10, 27, 'sp12_v_b_4')
// (10, 28, 'sp12_v_b_3')
// (10, 29, 'sp12_h_r_0')
// (10, 29, 'sp12_v_b_0')
// (10, 29, 'sp4_h_r_12')
// (10, 29, 'sp4_h_r_43')
// (11, 29, 'sp12_h_r_3')
// (11, 29, 'sp4_h_l_43')
// (11, 29, 'sp4_h_r_25')
// (11, 29, 'sp4_h_r_3')
// (12, 29, 'sp12_h_r_4')
// (12, 29, 'sp4_h_r_14')
// (12, 29, 'sp4_h_r_36')
// (13, 29, 'sp12_h_r_7')
// (13, 29, 'sp4_h_l_36')
// (13, 29, 'sp4_h_r_27')
// (14, 29, 'sp12_h_r_8')
// (14, 29, 'sp4_h_r_38')
// (15, 29, 'sp12_h_r_11')
// (15, 29, 'sp4_h_l_38')
// (16, 29, 'sp12_h_r_12')
// (17, 29, 'sp12_h_r_15')
// (18, 29, 'sp12_h_r_16')
// (19, 29, 'sp12_h_r_19')
// (20, 29, 'sp12_h_r_20')
// (21, 29, 'sp12_h_r_23')
// (22, 17, 'sp12_v_t_23')
// (22, 18, 'sp12_v_b_23')
// (22, 19, 'sp12_v_b_20')
// (22, 20, 'sp12_v_b_19')
// (22, 21, 'local_g3_0')
// (22, 21, 'lutff_5/in_0')
// (22, 21, 'sp12_v_b_16')
// (22, 22, 'sp12_v_b_15')
// (22, 23, 'sp12_v_b_12')
// (22, 24, 'sp12_v_b_11')
// (22, 25, 'sp12_v_b_8')
// (22, 26, 'sp12_v_b_7')
// (22, 27, 'sp12_v_b_4')
// (22, 28, 'sp12_v_b_3')
// (22, 29, 'sp12_h_l_23')
// (22, 29, 'sp12_h_r_0')
// (22, 29, 'sp12_v_b_0')
// (23, 29, 'sp12_h_r_3')
// (24, 14, 'sp4_r_v_b_38')
// (24, 15, 'sp4_r_v_b_27')
// (24, 16, 'sp4_r_v_b_14')
// (24, 17, 'sp4_r_v_b_3')
// (24, 18, 'sp4_r_v_b_38')
// (24, 19, 'sp4_r_v_b_27')
// (24, 20, 'sp4_r_v_b_14')
// (24, 21, 'sp4_r_v_b_3')
// (24, 22, 'sp4_r_v_b_38')
// (24, 23, 'sp4_r_v_b_27')
// (24, 24, 'sp4_r_v_b_14')
// (24, 25, 'sp4_r_v_b_3')
// (24, 26, 'sp4_r_v_b_43')
// (24, 27, 'sp4_r_v_b_30')
// (24, 28, 'sp4_r_v_b_19')
// (24, 29, 'sp12_h_r_4')
// (24, 29, 'sp4_r_v_b_6')
// (25, 13, 'sp4_v_t_38')
// (25, 14, 'sp4_v_b_38')
// (25, 15, 'local_g2_3')
// (25, 15, 'ram/RADDR_8')
// (25, 15, 'sp4_v_b_27')
// (25, 16, 'sp4_v_b_14')
// (25, 17, 'local_g1_0')
// (25, 17, 'ram/RADDR_8')
// (25, 17, 'sp4_h_r_0')
// (25, 17, 'sp4_h_r_3')
// (25, 17, 'sp4_v_b_3')
// (25, 17, 'sp4_v_t_38')
// (25, 18, 'sp4_v_b_38')
// (25, 19, 'local_g2_3')
// (25, 19, 'ram/RADDR_8')
// (25, 19, 'sp4_v_b_27')
// (25, 20, 'sp4_v_b_14')
// (25, 21, 'local_g1_0')
// (25, 21, 'ram/RADDR_8')
// (25, 21, 'sp4_h_r_0')
// (25, 21, 'sp4_h_r_3')
// (25, 21, 'sp4_v_b_3')
// (25, 21, 'sp4_v_t_38')
// (25, 22, 'sp4_v_b_38')
// (25, 23, 'local_g2_3')
// (25, 23, 'ram/RADDR_8')
// (25, 23, 'sp4_v_b_27')
// (25, 24, 'sp4_v_b_14')
// (25, 25, 'local_g0_3')
// (25, 25, 'ram/RADDR_8')
// (25, 25, 'sp4_h_r_3')
// (25, 25, 'sp4_v_b_3')
// (25, 25, 'sp4_v_t_43')
// (25, 26, 'sp4_v_b_43')
// (25, 27, 'local_g3_6')
// (25, 27, 'ram/RADDR_8')
// (25, 27, 'sp4_v_b_30')
// (25, 28, 'sp4_v_b_19')
// (25, 29, 'local_g0_1')
// (25, 29, 'ram/RADDR_8')
// (25, 29, 'sp12_h_r_7')
// (25, 29, 'sp4_h_r_1')
// (25, 29, 'sp4_v_b_6')
// (26, 17, 'sp4_h_r_13')
// (26, 17, 'sp4_h_r_14')
// (26, 21, 'local_g0_6')
// (26, 21, 'lutff_2/in_0')
// (26, 21, 'sp4_h_r_13')
// (26, 21, 'sp4_h_r_14')
// (26, 25, 'sp4_h_r_14')
// (26, 29, 'sp12_h_r_8')
// (26, 29, 'sp4_h_r_12')
// (27, 17, 'sp4_h_r_24')
// (27, 17, 'sp4_h_r_27')
// (27, 21, 'sp4_h_r_24')
// (27, 21, 'sp4_h_r_27')
// (27, 25, 'sp4_h_r_27')
// (27, 29, 'sp12_h_r_11')
// (27, 29, 'sp4_h_r_25')
// (28, 17, 'sp4_h_r_37')
// (28, 17, 'sp4_h_r_38')
// (28, 21, 'sp4_h_r_37')
// (28, 21, 'sp4_h_r_38')
// (28, 25, 'sp4_h_r_38')
// (28, 29, 'sp12_h_r_12')
// (28, 29, 'sp4_h_r_36')
// (29, 17, 'sp4_h_l_37')
// (29, 17, 'sp4_h_l_38')
// (29, 17, 'sp4_h_r_0')
// (29, 21, 'sp4_h_l_37')
// (29, 21, 'sp4_h_l_38')
// (29, 21, 'sp4_h_r_0')
// (29, 25, 'sp4_h_l_38')
// (29, 25, 'sp4_h_r_0')
// (29, 29, 'sp12_h_r_15')
// (29, 29, 'sp4_h_l_36')
// (29, 29, 'sp4_h_r_1')
// (30, 17, 'sp4_h_r_13')
// (30, 21, 'sp4_h_r_13')
// (30, 25, 'sp4_h_r_13')
// (30, 29, 'sp12_h_r_16')
// (30, 29, 'sp4_h_r_12')
// (31, 17, 'sp4_h_r_24')
// (31, 21, 'sp4_h_r_24')
// (31, 25, 'sp4_h_r_24')
// (31, 29, 'sp12_h_r_19')
// (31, 29, 'sp4_h_r_25')
// (32, 17, 'sp4_h_r_37')
// (32, 21, 'sp4_h_r_37')
// (32, 25, 'sp4_h_r_37')
// (32, 28, 'neigh_op_tnr_2')
// (32, 28, 'neigh_op_tnr_6')
// (32, 29, 'neigh_op_rgt_2')
// (32, 29, 'neigh_op_rgt_6')
// (32, 29, 'sp12_h_r_20')
// (32, 29, 'sp4_h_r_36')
// (32, 30, 'neigh_op_bnr_2')
// (32, 30, 'neigh_op_bnr_6')
// (33, 17, 'span4_horz_37')
// (33, 17, 'span4_vert_t_14')
// (33, 18, 'span4_vert_b_14')
// (33, 19, 'span4_vert_b_10')
// (33, 20, 'span4_vert_b_6')
// (33, 21, 'span4_horz_37')
// (33, 21, 'span4_vert_b_2')
// (33, 21, 'span4_vert_t_14')
// (33, 22, 'span4_vert_b_14')
// (33, 23, 'span4_vert_b_10')
// (33, 24, 'span4_vert_b_6')
// (33, 25, 'span4_horz_37')
// (33, 25, 'span4_vert_b_2')
// (33, 25, 'span4_vert_t_14')
// (33, 26, 'span4_vert_b_14')
// (33, 27, 'span4_vert_b_10')
// (33, 28, 'span4_vert_b_6')
// (33, 29, 'io_1/D_IN_0')
// (33, 29, 'io_1/PAD')
// (33, 29, 'span12_horz_20')
// (33, 29, 'span4_horz_36')
// (33, 29, 'span4_vert_b_2')

reg io_0_20_0 = 0;
// (0, 17, 'span4_vert_t_12')
// (0, 18, 'span4_vert_b_12')
// (0, 19, 'span4_vert_b_8')
// (0, 20, 'io_0/D_OUT_0')
// (0, 20, 'io_0/PAD')
// (0, 20, 'local_g0_4')
// (0, 20, 'span4_vert_b_4')
// (0, 21, 'span4_horz_1')
// (0, 21, 'span4_vert_b_0')
// (1, 21, 'sp4_h_r_12')
// (2, 21, 'sp4_h_r_25')
// (3, 21, 'sp4_h_r_36')
// (4, 21, 'sp4_h_l_36')
// (4, 21, 'sp4_h_r_5')
// (5, 21, 'sp4_h_r_16')
// (6, 20, 'neigh_op_tnr_4')
// (6, 21, 'neigh_op_rgt_4')
// (6, 21, 'sp4_h_r_29')
// (6, 22, 'neigh_op_bnr_4')
// (7, 20, 'neigh_op_top_4')
// (7, 21, 'lutff_4/out')
// (7, 21, 'sp4_h_r_40')
// (7, 22, 'neigh_op_bot_4')
// (8, 20, 'neigh_op_tnl_4')
// (8, 21, 'neigh_op_lft_4')
// (8, 21, 'sp4_h_l_40')
// (8, 22, 'neigh_op_bnl_4')

reg io_0_20_1 = 0;
// (0, 17, 'span4_vert_t_15')
// (0, 18, 'span4_vert_b_15')
// (0, 19, 'span4_vert_b_11')
// (0, 20, 'io_1/D_OUT_0')
// (0, 20, 'io_1/PAD')
// (0, 20, 'local_g0_7')
// (0, 20, 'span4_vert_b_7')
// (0, 21, 'span4_horz_43')
// (0, 21, 'span4_vert_b_3')
// (1, 21, 'sp4_h_l_43')
// (1, 21, 'sp4_h_r_10')
// (2, 21, 'sp4_h_r_23')
// (3, 21, 'sp4_h_r_34')
// (4, 21, 'sp4_h_r_47')
// (5, 21, 'sp4_h_l_47')
// (5, 21, 'sp4_h_r_10')
// (6, 20, 'neigh_op_tnr_1')
// (6, 21, 'neigh_op_rgt_1')
// (6, 21, 'sp4_h_r_23')
// (6, 22, 'neigh_op_bnr_1')
// (7, 20, 'neigh_op_top_1')
// (7, 21, 'lutff_1/out')
// (7, 21, 'sp4_h_r_34')
// (7, 22, 'neigh_op_bot_1')
// (8, 20, 'neigh_op_tnl_1')
// (8, 21, 'neigh_op_lft_1')
// (8, 21, 'sp4_h_r_47')
// (8, 22, 'neigh_op_bnl_1')
// (9, 21, 'sp4_h_l_47')

reg io_0_18_0 = 0;
// (0, 18, 'io_0/D_OUT_0')
// (0, 18, 'io_0/PAD')
// (0, 18, 'local_g1_3')
// (0, 18, 'span4_horz_19')
// (1, 18, 'sp4_h_r_30')
// (2, 18, 'sp4_h_r_43')
// (3, 18, 'sp4_h_l_43')
// (3, 18, 'sp4_h_r_3')
// (4, 18, 'sp4_h_r_14')
// (5, 18, 'sp4_h_r_27')
// (6, 18, 'sp4_h_r_38')
// (6, 19, 'sp4_r_v_b_38')
// (6, 20, 'neigh_op_tnr_7')
// (6, 20, 'sp4_r_v_b_27')
// (6, 21, 'neigh_op_rgt_7')
// (6, 21, 'sp4_r_v_b_14')
// (6, 22, 'neigh_op_bnr_7')
// (6, 22, 'sp4_r_v_b_3')
// (7, 18, 'sp4_h_l_38')
// (7, 18, 'sp4_v_t_38')
// (7, 19, 'sp4_v_b_38')
// (7, 20, 'neigh_op_top_7')
// (7, 20, 'sp4_v_b_27')
// (7, 21, 'lutff_7/out')
// (7, 21, 'sp4_v_b_14')
// (7, 22, 'neigh_op_bot_7')
// (7, 22, 'sp4_v_b_3')
// (8, 20, 'neigh_op_tnl_7')
// (8, 21, 'neigh_op_lft_7')
// (8, 22, 'neigh_op_bnl_7')

wire io_33_31_0;
// (0, 19, 'span12_horz_0')
// (1, 19, 'sp12_h_r_3')
// (2, 19, 'sp12_h_r_4')
// (3, 19, 'sp12_h_r_7')
// (4, 19, 'sp12_h_r_8')
// (5, 19, 'sp12_h_r_11')
// (6, 19, 'sp12_h_r_12')
// (7, 19, 'sp12_h_r_15')
// (8, 15, 'local_g1_1')
// (8, 15, 'ram/RADDR_7')
// (8, 15, 'sp4_h_r_9')
// (8, 17, 'local_g0_2')
// (8, 17, 'ram/RADDR_7')
// (8, 17, 'sp4_h_r_10')
// (8, 19, 'local_g0_0')
// (8, 19, 'ram/RADDR_7')
// (8, 19, 'sp12_h_r_16')
// (8, 21, 'local_g0_2')
// (8, 21, 'ram/RADDR_7')
// (8, 21, 'sp4_h_r_10')
// (8, 23, 'local_g1_1')
// (8, 23, 'ram/RADDR_7')
// (8, 23, 'sp4_h_r_1')
// (8, 25, 'local_g0_6')
// (8, 25, 'ram/RADDR_7')
// (8, 25, 'sp4_h_r_6')
// (8, 27, 'local_g1_1')
// (8, 27, 'ram/RADDR_7')
// (8, 27, 'sp4_h_r_9')
// (8, 29, 'local_g0_2')
// (8, 29, 'ram/RADDR_7')
// (8, 29, 'sp4_h_r_2')
// (9, 15, 'sp4_h_r_20')
// (9, 17, 'sp4_h_r_23')
// (9, 19, 'sp12_h_r_19')
// (9, 21, 'sp4_h_r_23')
// (9, 23, 'sp4_h_r_12')
// (9, 25, 'sp4_h_r_19')
// (9, 27, 'sp4_h_r_20')
// (9, 29, 'sp4_h_r_15')
// (10, 15, 'sp4_h_r_33')
// (10, 17, 'sp4_h_r_34')
// (10, 19, 'sp12_h_r_20')
// (10, 21, 'sp4_h_r_34')
// (10, 23, 'sp4_h_r_25')
// (10, 25, 'sp4_h_r_30')
// (10, 27, 'sp4_h_r_33')
// (10, 29, 'sp4_h_r_26')
// (11, 12, 'sp4_r_v_b_41')
// (11, 13, 'sp4_r_v_b_28')
// (11, 14, 'sp4_r_v_b_17')
// (11, 15, 'sp4_h_r_44')
// (11, 15, 'sp4_r_v_b_4')
// (11, 17, 'sp4_h_r_47')
// (11, 18, 'sp4_r_v_b_47')
// (11, 19, 'sp12_h_r_23')
// (11, 19, 'sp4_r_v_b_34')
// (11, 20, 'sp4_r_v_b_23')
// (11, 20, 'sp4_r_v_b_45')
// (11, 21, 'sp4_h_r_47')
// (11, 21, 'sp4_r_v_b_10')
// (11, 21, 'sp4_r_v_b_32')
// (11, 22, 'sp4_r_v_b_21')
// (11, 22, 'sp4_r_v_b_43')
// (11, 23, 'sp4_h_r_36')
// (11, 23, 'sp4_r_v_b_30')
// (11, 23, 'sp4_r_v_b_8')
// (11, 24, 'sp4_r_v_b_19')
// (11, 24, 'sp4_r_v_b_41')
// (11, 25, 'sp4_h_r_43')
// (11, 25, 'sp4_r_v_b_28')
// (11, 25, 'sp4_r_v_b_6')
// (11, 26, 'sp4_r_v_b_17')
// (11, 26, 'sp4_r_v_b_39')
// (11, 27, 'sp4_h_r_44')
// (11, 27, 'sp4_r_v_b_26')
// (11, 27, 'sp4_r_v_b_4')
// (11, 28, 'sp4_r_v_b_15')
// (11, 29, 'sp4_h_r_39')
// (11, 29, 'sp4_r_v_b_2')
// (12, 7, 'sp12_v_t_23')
// (12, 8, 'sp12_v_b_23')
// (12, 9, 'sp12_v_b_20')
// (12, 10, 'sp12_v_b_19')
// (12, 11, 'sp12_v_b_16')
// (12, 11, 'sp4_v_t_41')
// (12, 12, 'sp12_v_b_15')
// (12, 12, 'sp4_v_b_41')
// (12, 13, 'sp12_v_b_12')
// (12, 13, 'sp4_v_b_28')
// (12, 14, 'sp12_v_b_11')
// (12, 14, 'sp4_v_b_17')
// (12, 15, 'sp12_v_b_8')
// (12, 15, 'sp4_h_l_44')
// (12, 15, 'sp4_v_b_4')
// (12, 16, 'sp12_v_b_7')
// (12, 17, 'sp12_v_b_4')
// (12, 17, 'sp4_h_l_47')
// (12, 17, 'sp4_v_t_47')
// (12, 18, 'sp12_v_b_3')
// (12, 18, 'sp4_v_b_47')
// (12, 19, 'sp12_h_l_23')
// (12, 19, 'sp12_h_r_0')
// (12, 19, 'sp12_v_b_0')
// (12, 19, 'sp12_v_t_23')
// (12, 19, 'sp4_v_b_34')
// (12, 19, 'sp4_v_t_45')
// (12, 20, 'sp12_v_b_23')
// (12, 20, 'sp4_v_b_23')
// (12, 20, 'sp4_v_b_45')
// (12, 21, 'sp12_v_b_20')
// (12, 21, 'sp4_h_l_47')
// (12, 21, 'sp4_v_b_10')
// (12, 21, 'sp4_v_b_32')
// (12, 21, 'sp4_v_t_43')
// (12, 22, 'sp12_v_b_19')
// (12, 22, 'sp4_v_b_21')
// (12, 22, 'sp4_v_b_43')
// (12, 23, 'sp12_v_b_16')
// (12, 23, 'sp4_h_l_36')
// (12, 23, 'sp4_v_b_30')
// (12, 23, 'sp4_v_b_8')
// (12, 23, 'sp4_v_t_41')
// (12, 24, 'sp12_v_b_15')
// (12, 24, 'sp4_v_b_19')
// (12, 24, 'sp4_v_b_41')
// (12, 25, 'sp12_v_b_12')
// (12, 25, 'sp4_h_l_43')
// (12, 25, 'sp4_v_b_28')
// (12, 25, 'sp4_v_b_6')
// (12, 25, 'sp4_v_t_39')
// (12, 26, 'sp12_v_b_11')
// (12, 26, 'sp4_v_b_17')
// (12, 26, 'sp4_v_b_39')
// (12, 27, 'sp12_v_b_8')
// (12, 27, 'sp4_h_l_44')
// (12, 27, 'sp4_v_b_26')
// (12, 27, 'sp4_v_b_4')
// (12, 28, 'sp12_v_b_7')
// (12, 28, 'sp4_v_b_15')
// (12, 29, 'sp12_v_b_4')
// (12, 29, 'sp4_h_l_39')
// (12, 29, 'sp4_v_b_2')
// (12, 30, 'sp12_v_b_3')
// (12, 31, 'sp12_h_r_0')
// (12, 31, 'sp12_v_b_0')
// (13, 19, 'sp12_h_r_3')
// (13, 31, 'sp12_h_r_3')
// (14, 19, 'sp12_h_r_4')
// (14, 31, 'sp12_h_r_4')
// (15, 19, 'sp12_h_r_7')
// (15, 31, 'sp12_h_r_7')
// (16, 19, 'sp12_h_r_8')
// (16, 31, 'sp12_h_r_8')
// (17, 19, 'sp12_h_r_11')
// (17, 31, 'sp12_h_r_11')
// (18, 19, 'sp12_h_r_12')
// (18, 31, 'sp12_h_r_12')
// (19, 19, 'sp12_h_r_15')
// (19, 31, 'sp12_h_r_15')
// (20, 19, 'local_g1_0')
// (20, 19, 'lutff_5/in_2')
// (20, 19, 'sp12_h_r_16')
// (20, 31, 'sp12_h_r_16')
// (21, 19, 'sp12_h_r_19')
// (21, 31, 'sp12_h_r_19')
// (22, 19, 'sp12_h_r_20')
// (22, 31, 'sp12_h_r_20')
// (23, 16, 'sp4_r_v_b_46')
// (23, 17, 'sp4_r_v_b_35')
// (23, 18, 'sp4_r_v_b_22')
// (23, 18, 'sp4_r_v_b_47')
// (23, 19, 'sp12_h_r_23')
// (23, 19, 'sp4_r_v_b_11')
// (23, 19, 'sp4_r_v_b_34')
// (23, 20, 'sp4_r_v_b_23')
// (23, 20, 'sp4_r_v_b_45')
// (23, 21, 'local_g2_2')
// (23, 21, 'lutff_0/in_2')
// (23, 21, 'sp4_r_v_b_10')
// (23, 21, 'sp4_r_v_b_32')
// (23, 22, 'sp4_r_v_b_21')
// (23, 23, 'sp4_r_v_b_8')
// (23, 31, 'sp12_h_r_23')
// (24, 15, 'sp4_h_r_11')
// (24, 15, 'sp4_v_t_46')
// (24, 16, 'sp4_v_b_46')
// (24, 17, 'sp4_h_r_10')
// (24, 17, 'sp4_v_b_35')
// (24, 17, 'sp4_v_t_47')
// (24, 18, 'sp4_v_b_22')
// (24, 18, 'sp4_v_b_47')
// (24, 19, 'sp12_h_l_23')
// (24, 19, 'sp12_h_r_0')
// (24, 19, 'sp12_v_t_23')
// (24, 19, 'sp4_v_b_11')
// (24, 19, 'sp4_v_b_34')
// (24, 19, 'sp4_v_t_45')
// (24, 20, 'sp12_v_b_23')
// (24, 20, 'sp4_v_b_23')
// (24, 20, 'sp4_v_b_45')
// (24, 21, 'sp12_v_b_20')
// (24, 21, 'sp4_h_r_4')
// (24, 21, 'sp4_v_b_10')
// (24, 21, 'sp4_v_b_32')
// (24, 22, 'sp12_v_b_19')
// (24, 22, 'sp4_v_b_21')
// (24, 23, 'sp12_v_b_16')
// (24, 23, 'sp4_h_r_7')
// (24, 23, 'sp4_v_b_8')
// (24, 24, 'sp12_v_b_15')
// (24, 25, 'sp12_v_b_12')
// (24, 26, 'sp12_v_b_11')
// (24, 27, 'sp12_v_b_8')
// (24, 28, 'sp12_v_b_7')
// (24, 28, 'sp4_r_v_b_45')
// (24, 29, 'sp12_v_b_4')
// (24, 29, 'sp4_r_v_b_32')
// (24, 30, 'sp12_v_b_3')
// (24, 30, 'sp4_r_v_b_21')
// (24, 31, 'sp12_h_l_23')
// (24, 31, 'sp12_h_r_0')
// (24, 31, 'sp12_v_b_0')
// (24, 31, 'sp4_r_v_b_8')
// (25, 15, 'local_g0_6')
// (25, 15, 'ram/RADDR_7')
// (25, 15, 'sp4_h_r_22')
// (25, 17, 'local_g1_7')
// (25, 17, 'ram/RADDR_7')
// (25, 17, 'sp4_h_r_23')
// (25, 19, 'local_g1_3')
// (25, 19, 'ram/RADDR_7')
// (25, 19, 'sp12_h_r_3')
// (25, 21, 'local_g1_1')
// (25, 21, 'ram/RADDR_7')
// (25, 21, 'sp4_h_r_17')
// (25, 23, 'local_g0_2')
// (25, 23, 'ram/RADDR_7')
// (25, 23, 'sp4_h_r_18')
// (25, 24, 'sp4_r_v_b_36')
// (25, 24, 'sp4_r_v_b_41')
// (25, 25, 'local_g0_4')
// (25, 25, 'ram/RADDR_7')
// (25, 25, 'sp4_r_v_b_25')
// (25, 25, 'sp4_r_v_b_28')
// (25, 26, 'sp4_r_v_b_12')
// (25, 26, 'sp4_r_v_b_17')
// (25, 27, 'local_g1_1')
// (25, 27, 'ram/RADDR_7')
// (25, 27, 'sp4_r_v_b_1')
// (25, 27, 'sp4_r_v_b_4')
// (25, 27, 'sp4_v_t_45')
// (25, 28, 'sp4_v_b_45')
// (25, 29, 'local_g2_0')
// (25, 29, 'ram/RADDR_7')
// (25, 29, 'sp4_v_b_32')
// (25, 30, 'sp4_v_b_21')
// (25, 31, 'sp12_h_r_3')
// (25, 31, 'sp4_h_r_8')
// (25, 31, 'sp4_v_b_8')
// (26, 15, 'sp4_h_r_35')
// (26, 17, 'sp4_h_r_34')
// (26, 19, 'sp12_h_r_4')
// (26, 21, 'sp4_h_r_28')
// (26, 23, 'sp4_h_r_31')
// (26, 23, 'sp4_v_t_36')
// (26, 23, 'sp4_v_t_41')
// (26, 24, 'sp4_v_b_36')
// (26, 24, 'sp4_v_b_41')
// (26, 25, 'sp4_v_b_25')
// (26, 25, 'sp4_v_b_28')
// (26, 26, 'sp4_v_b_12')
// (26, 26, 'sp4_v_b_17')
// (26, 27, 'sp4_h_r_1')
// (26, 27, 'sp4_h_r_4')
// (26, 27, 'sp4_v_b_1')
// (26, 27, 'sp4_v_b_4')
// (26, 31, 'sp12_h_r_4')
// (26, 31, 'sp4_h_r_21')
// (27, 15, 'sp4_h_r_46')
// (27, 17, 'sp4_h_r_47')
// (27, 19, 'sp12_h_r_7')
// (27, 21, 'sp4_h_r_41')
// (27, 23, 'sp4_h_r_42')
// (27, 27, 'sp4_h_r_12')
// (27, 27, 'sp4_h_r_17')
// (27, 31, 'sp12_h_r_7')
// (27, 31, 'sp4_h_r_32')
// (28, 15, 'sp4_h_l_46')
// (28, 17, 'sp4_h_l_47')
// (28, 19, 'sp12_h_r_8')
// (28, 21, 'sp4_h_l_41')
// (28, 23, 'sp4_h_l_42')
// (28, 23, 'sp4_h_r_4')
// (28, 27, 'sp4_h_r_25')
// (28, 27, 'sp4_h_r_28')
// (28, 31, 'sp12_h_r_8')
// (28, 31, 'sp4_h_r_45')
// (29, 19, 'sp12_h_r_11')
// (29, 23, 'sp4_h_r_17')
// (29, 27, 'sp4_h_r_36')
// (29, 27, 'sp4_h_r_41')
// (29, 31, 'sp12_h_r_11')
// (29, 31, 'sp4_h_l_45')
// (29, 31, 'sp4_h_r_5')
// (30, 19, 'sp12_h_r_12')
// (30, 23, 'sp4_h_r_28')
// (30, 27, 'sp4_h_l_36')
// (30, 27, 'sp4_h_l_41')
// (30, 27, 'sp4_h_r_1')
// (30, 31, 'sp12_h_r_12')
// (30, 31, 'sp4_h_r_16')
// (31, 19, 'sp12_h_r_15')
// (31, 23, 'sp4_h_r_41')
// (31, 27, 'sp4_h_r_12')
// (31, 31, 'sp12_h_r_15')
// (31, 31, 'sp4_h_r_29')
// (32, 19, 'sp12_h_r_16')
// (32, 23, 'sp4_h_l_41')
// (32, 23, 'sp4_h_r_1')
// (32, 27, 'sp4_h_r_25')
// (32, 30, 'neigh_op_tnr_0')
// (32, 30, 'neigh_op_tnr_4')
// (32, 31, 'neigh_op_rgt_0')
// (32, 31, 'neigh_op_rgt_4')
// (32, 31, 'sp12_h_r_16')
// (32, 31, 'sp4_h_r_40')
// (32, 32, 'neigh_op_bnr_0')
// (32, 32, 'neigh_op_bnr_4')
// (33, 19, 'span12_horz_16')
// (33, 23, 'span4_horz_1')
// (33, 23, 'span4_vert_t_12')
// (33, 24, 'span4_vert_b_12')
// (33, 25, 'span4_vert_b_8')
// (33, 26, 'span4_vert_b_4')
// (33, 27, 'span4_horz_25')
// (33, 27, 'span4_vert_b_0')
// (33, 27, 'span4_vert_t_12')
// (33, 28, 'span4_vert_b_12')
// (33, 29, 'span4_vert_b_8')
// (33, 30, 'span4_vert_b_4')
// (33, 31, 'io_0/D_IN_0')
// (33, 31, 'io_0/PAD')
// (33, 31, 'span12_horz_16')
// (33, 31, 'span4_horz_40')
// (33, 31, 'span4_vert_b_0')

reg io_0_22_0 = 0;
// (0, 22, 'io_0/D_OUT_0')
// (0, 22, 'io_0/PAD')
// (0, 22, 'local_g1_5')
// (0, 22, 'span12_horz_5')
// (1, 22, 'sp12_h_r_6')
// (2, 22, 'sp12_h_r_9')
// (3, 22, 'sp12_h_r_10')
// (4, 22, 'sp12_h_r_13')
// (5, 22, 'sp12_h_r_14')
// (6, 21, 'neigh_op_tnr_5')
// (6, 22, 'neigh_op_rgt_5')
// (6, 22, 'sp12_h_r_17')
// (6, 23, 'neigh_op_bnr_5')
// (7, 21, 'neigh_op_top_5')
// (7, 22, 'lutff_5/out')
// (7, 22, 'sp12_h_r_18')
// (7, 23, 'neigh_op_bot_5')
// (8, 21, 'neigh_op_tnl_5')
// (8, 22, 'neigh_op_lft_5')
// (8, 22, 'sp12_h_r_21')
// (8, 23, 'neigh_op_bnl_5')
// (9, 22, 'sp12_h_r_22')
// (10, 22, 'sp12_h_l_22')

reg io_0_22_1 = 0;
// (0, 22, 'io_1/D_OUT_0')
// (0, 22, 'io_1/PAD')
// (0, 22, 'local_g0_1')
// (0, 22, 'span4_horz_41')
// (1, 22, 'sp4_h_l_41')
// (1, 22, 'sp4_h_r_1')
// (2, 22, 'sp4_h_r_12')
// (3, 22, 'sp4_h_r_25')
// (4, 22, 'sp4_h_r_36')
// (5, 22, 'sp4_h_l_36')
// (5, 22, 'sp4_h_r_10')
// (6, 21, 'neigh_op_tnr_1')
// (6, 22, 'neigh_op_rgt_1')
// (6, 22, 'sp4_h_r_23')
// (6, 23, 'neigh_op_bnr_1')
// (7, 21, 'neigh_op_top_1')
// (7, 22, 'lutff_1/out')
// (7, 22, 'sp4_h_r_34')
// (7, 23, 'neigh_op_bot_1')
// (8, 21, 'neigh_op_tnl_1')
// (8, 22, 'neigh_op_lft_1')
// (8, 22, 'sp4_h_r_47')
// (8, 23, 'neigh_op_bnl_1')
// (9, 22, 'sp4_h_l_47')

wire n18;
// (0, 22, 'logic_op_tnr_0')
// (0, 23, 'logic_op_rgt_0')
// (0, 23, 'span4_horz_5')
// (0, 24, 'logic_op_bnr_0')
// (1, 20, 'sp4_r_v_b_36')
// (1, 21, 'sp4_r_v_b_25')
// (1, 21, 'sp4_r_v_b_41')
// (1, 22, 'neigh_op_top_0')
// (1, 22, 'sp4_r_v_b_12')
// (1, 22, 'sp4_r_v_b_28')
// (1, 22, 'sp4_r_v_b_44')
// (1, 23, 'lutff_0/out')
// (1, 23, 'sp4_h_r_16')
// (1, 23, 'sp4_r_v_b_1')
// (1, 23, 'sp4_r_v_b_17')
// (1, 23, 'sp4_r_v_b_33')
// (1, 24, 'neigh_op_bot_0')
// (1, 24, 'sp4_r_v_b_20')
// (1, 24, 'sp4_r_v_b_4')
// (1, 25, 'sp4_r_v_b_9')
// (2, 19, 'sp4_h_r_1')
// (2, 19, 'sp4_v_t_36')
// (2, 20, 'sp4_h_r_4')
// (2, 20, 'sp4_v_b_36')
// (2, 20, 'sp4_v_t_41')
// (2, 21, 'sp4_h_r_9')
// (2, 21, 'sp4_v_b_25')
// (2, 21, 'sp4_v_b_41')
// (2, 21, 'sp4_v_t_44')
// (2, 22, 'neigh_op_tnl_0')
// (2, 22, 'sp4_v_b_12')
// (2, 22, 'sp4_v_b_28')
// (2, 22, 'sp4_v_b_44')
// (2, 23, 'neigh_op_lft_0')
// (2, 23, 'sp4_h_r_29')
// (2, 23, 'sp4_v_b_1')
// (2, 23, 'sp4_v_b_17')
// (2, 23, 'sp4_v_b_33')
// (2, 24, 'neigh_op_bnl_0')
// (2, 24, 'sp4_v_b_20')
// (2, 24, 'sp4_v_b_4')
// (2, 25, 'sp4_v_b_9')
// (3, 19, 'sp4_h_r_12')
// (3, 20, 'sp4_h_r_17')
// (3, 21, 'sp4_h_r_20')
// (3, 23, 'sp4_h_r_40')
// (4, 19, 'sp4_h_r_25')
// (4, 20, 'sp4_h_r_28')
// (4, 21, 'sp4_h_r_33')
// (4, 23, 'sp4_h_l_40')
// (4, 23, 'sp4_h_r_8')
// (5, 17, 'sp4_r_v_b_47')
// (5, 18, 'sp4_r_v_b_34')
// (5, 19, 'sp4_h_r_36')
// (5, 19, 'sp4_r_v_b_23')
// (5, 20, 'sp4_h_r_41')
// (5, 20, 'sp4_r_v_b_10')
// (5, 21, 'sp4_h_r_44')
// (5, 23, 'sp4_h_r_21')
// (6, 16, 'sp4_v_t_47')
// (6, 17, 'sp4_v_b_47')
// (6, 18, 'sp4_v_b_34')
// (6, 19, 'sp4_h_l_36')
// (6, 19, 'sp4_h_r_4')
// (6, 19, 'sp4_v_b_23')
// (6, 20, 'local_g0_2')
// (6, 20, 'lutff_global/cen')
// (6, 20, 'sp4_h_l_41')
// (6, 20, 'sp4_h_r_7')
// (6, 20, 'sp4_v_b_10')
// (6, 21, 'local_g1_0')
// (6, 21, 'lutff_2/in_3')
// (6, 21, 'sp4_h_l_44')
// (6, 21, 'sp4_h_r_0')
// (6, 21, 'sp4_h_r_5')
// (6, 23, 'sp4_h_r_32')
// (7, 19, 'local_g1_1')
// (7, 19, 'lutff_0/in_2')
// (7, 19, 'lutff_3/in_1')
// (7, 19, 'sp4_h_r_17')
// (7, 20, 'local_g0_2')
// (7, 20, 'lutff_global/cen')
// (7, 20, 'sp4_h_r_18')
// (7, 20, 'sp4_r_v_b_39')
// (7, 21, 'local_g0_0')
// (7, 21, 'local_g1_0')
// (7, 21, 'lutff_1/in_0')
// (7, 21, 'lutff_4/in_2')
// (7, 21, 'lutff_5/in_2')
// (7, 21, 'lutff_7/in_0')
// (7, 21, 'sp4_h_r_13')
// (7, 21, 'sp4_h_r_16')
// (7, 21, 'sp4_r_v_b_26')
// (7, 22, 'local_g2_7')
// (7, 22, 'lutff_1/in_2')
// (7, 22, 'lutff_5/in_0')
// (7, 22, 'sp4_r_v_b_15')
// (7, 23, 'sp4_h_r_45')
// (7, 23, 'sp4_r_v_b_2')
// (8, 19, 'sp4_h_r_28')
// (8, 19, 'sp4_v_t_39')
// (8, 20, 'sp4_h_r_31')
// (8, 20, 'sp4_v_b_39')
// (8, 21, 'sp4_h_r_24')
// (8, 21, 'sp4_h_r_29')
// (8, 21, 'sp4_v_b_26')
// (8, 22, 'sp4_v_b_15')
// (8, 23, 'sp4_h_l_45')
// (8, 23, 'sp4_v_b_2')
// (9, 19, 'sp4_h_r_41')
// (9, 20, 'sp4_h_r_42')
// (9, 21, 'sp4_h_r_37')
// (9, 21, 'sp4_h_r_40')
// (10, 19, 'sp4_h_l_41')
// (10, 20, 'sp4_h_l_42')
// (10, 21, 'sp4_h_l_37')
// (10, 21, 'sp4_h_l_40')

wire io_0_27_0;
// (0, 23, 'span4_horz_25')
// (0, 23, 'span4_vert_t_12')
// (0, 24, 'span4_vert_b_12')
// (0, 25, 'span4_vert_b_8')
// (0, 26, 'span4_vert_b_4')
// (0, 27, 'io_0/D_IN_0')
// (0, 27, 'io_0/PAD')
// (0, 27, 'span12_horz_0')
// (0, 27, 'span4_vert_b_0')
// (1, 23, 'local_g2_4')
// (1, 23, 'lutff_0/in_2')
// (1, 23, 'sp4_h_r_36')
// (1, 26, 'neigh_op_tnl_0')
// (1, 26, 'neigh_op_tnl_4')
// (1, 27, 'neigh_op_lft_0')
// (1, 27, 'neigh_op_lft_4')
// (1, 27, 'sp12_h_r_3')
// (1, 28, 'neigh_op_bnl_0')
// (1, 28, 'neigh_op_bnl_4')
// (2, 23, 'sp4_h_l_36')
// (2, 27, 'sp12_h_r_4')
// (3, 27, 'sp12_h_r_7')
// (4, 27, 'sp12_h_r_8')
// (5, 27, 'sp12_h_r_11')
// (6, 27, 'sp12_h_r_12')
// (7, 27, 'sp12_h_r_15')
// (8, 27, 'sp12_h_r_16')
// (9, 27, 'sp12_h_r_19')
// (9, 27, 'sp4_h_r_11')
// (10, 27, 'sp12_h_r_20')
// (10, 27, 'sp4_h_r_22')
// (11, 27, 'sp12_h_r_23')
// (11, 27, 'sp4_h_r_35')
// (12, 27, 'sp12_h_l_23')
// (12, 27, 'sp4_h_r_46')
// (13, 27, 'sp4_h_l_46')
// (13, 27, 'sp4_h_r_7')
// (14, 27, 'sp4_h_r_18')
// (15, 27, 'sp4_h_r_31')
// (16, 20, 'sp4_r_v_b_44')
// (16, 21, 'sp4_r_v_b_33')
// (16, 22, 'sp4_r_v_b_20')
// (16, 23, 'sp4_r_v_b_9')
// (16, 24, 'sp4_r_v_b_36')
// (16, 25, 'sp4_r_v_b_25')
// (16, 26, 'sp4_r_v_b_12')
// (16, 27, 'sp4_h_r_42')
// (16, 27, 'sp4_r_v_b_1')
// (17, 19, 'sp4_v_t_44')
// (17, 20, 'sp4_v_b_44')
// (17, 21, 'local_g2_1')
// (17, 21, 'lutff_4/in_3')
// (17, 21, 'sp4_v_b_33')
// (17, 22, 'sp4_v_b_20')
// (17, 23, 'sp4_v_b_9')
// (17, 23, 'sp4_v_t_36')
// (17, 24, 'sp4_v_b_36')
// (17, 25, 'sp4_v_b_25')
// (17, 26, 'sp4_v_b_12')
// (17, 27, 'sp4_h_l_42')
// (17, 27, 'sp4_v_b_1')

wire io_0_25_0;
// (0, 25, 'io_0/D_IN_0')
// (0, 25, 'io_0/PAD')
// (0, 25, 'span4_horz_40')
// (1, 21, 'sp4_v_t_46')
// (1, 22, 'sp4_v_b_46')
// (1, 23, 'local_g3_3')
// (1, 23, 'lutff_0/in_0')
// (1, 23, 'sp4_v_b_35')
// (1, 24, 'neigh_op_tnl_0')
// (1, 24, 'neigh_op_tnl_4')
// (1, 24, 'sp4_v_b_22')
// (1, 25, 'neigh_op_lft_0')
// (1, 25, 'neigh_op_lft_4')
// (1, 25, 'sp4_h_l_40')
// (1, 25, 'sp4_v_b_11')
// (1, 26, 'neigh_op_bnl_0')
// (1, 26, 'neigh_op_bnl_4')

wire n21;
// (1, 21, 'sp12_h_r_1')
// (2, 21, 'sp12_h_r_2')
// (3, 21, 'sp12_h_r_5')
// (4, 21, 'sp12_h_r_6')
// (5, 21, 'sp12_h_r_9')
// (6, 21, 'sp12_h_r_10')
// (7, 21, 'local_g0_5')
// (7, 21, 'lutff_4/in_1')
// (7, 21, 'sp12_h_r_13')
// (8, 21, 'sp12_h_r_14')
// (9, 21, 'sp12_h_r_17')
// (10, 21, 'sp12_h_r_18')
// (11, 21, 'sp12_h_r_21')
// (12, 21, 'sp12_h_r_22')
// (13, 21, 'sp12_h_l_22')
// (13, 21, 'sp12_h_r_1')
// (14, 21, 'sp12_h_r_2')
// (15, 21, 'sp12_h_r_5')
// (16, 21, 'sp12_h_r_6')
// (17, 21, 'sp12_h_r_9')
// (18, 21, 'sp12_h_r_10')
// (19, 21, 'sp12_h_r_13')
// (20, 21, 'sp12_h_r_14')
// (21, 21, 'sp12_h_r_17')
// (22, 21, 'sp12_h_r_18')
// (23, 20, 'neigh_op_tnr_7')
// (23, 21, 'neigh_op_rgt_7')
// (23, 21, 'sp12_h_r_21')
// (23, 22, 'neigh_op_bnr_7')
// (24, 20, 'neigh_op_top_7')
// (24, 21, 'lutff_7/out')
// (24, 21, 'sp12_h_r_22')
// (24, 22, 'neigh_op_bot_7')
// (25, 20, 'neigh_op_tnl_7')
// (25, 21, 'neigh_op_lft_7')
// (25, 21, 'sp12_h_l_22')
// (25, 22, 'neigh_op_bnl_7')

wire n22;
// (1, 22, 'sp12_h_r_1')
// (2, 22, 'sp12_h_r_2')
// (3, 22, 'sp12_h_r_5')
// (4, 22, 'sp12_h_r_6')
// (5, 22, 'sp12_h_r_9')
// (6, 22, 'sp12_h_r_10')
// (7, 22, 'local_g1_5')
// (7, 22, 'lutff_5/in_1')
// (7, 22, 'sp12_h_r_13')
// (8, 22, 'sp12_h_r_14')
// (9, 22, 'sp12_h_r_17')
// (10, 22, 'sp12_h_r_18')
// (11, 22, 'sp12_h_r_21')
// (12, 22, 'sp12_h_r_22')
// (13, 22, 'sp12_h_l_22')
// (13, 22, 'sp12_h_r_1')
// (14, 22, 'sp12_h_r_2')
// (15, 22, 'sp12_h_r_5')
// (16, 22, 'sp12_h_r_6')
// (17, 22, 'sp12_h_r_9')
// (18, 22, 'sp12_h_r_10')
// (19, 22, 'sp12_h_r_13')
// (20, 22, 'sp12_h_r_14')
// (21, 22, 'sp12_h_r_17')
// (22, 22, 'sp12_h_r_18')
// (23, 21, 'neigh_op_tnr_7')
// (23, 22, 'neigh_op_rgt_7')
// (23, 22, 'sp12_h_r_21')
// (23, 23, 'neigh_op_bnr_7')
// (24, 21, 'neigh_op_top_7')
// (24, 22, 'lutff_7/out')
// (24, 22, 'sp12_h_r_22')
// (24, 23, 'neigh_op_bot_7')
// (25, 21, 'neigh_op_tnl_7')
// (25, 22, 'neigh_op_lft_7')
// (25, 22, 'sp12_h_l_22')
// (25, 23, 'neigh_op_bnl_7')

wire io_3_33_1;
// (2, 18, 'sp4_r_v_b_47')
// (2, 19, 'sp4_r_v_b_34')
// (2, 20, 'sp4_r_v_b_23')
// (2, 20, 'sp4_r_v_b_41')
// (2, 21, 'sp4_r_v_b_10')
// (2, 21, 'sp4_r_v_b_28')
// (2, 22, 'sp4_r_v_b_17')
// (2, 22, 'sp4_r_v_b_47')
// (2, 23, 'sp4_r_v_b_34')
// (2, 23, 'sp4_r_v_b_4')
// (2, 24, 'sp4_r_v_b_23')
// (2, 24, 'sp4_r_v_b_45')
// (2, 25, 'sp4_r_v_b_10')
// (2, 25, 'sp4_r_v_b_32')
// (2, 26, 'sp4_r_v_b_21')
// (2, 27, 'sp4_r_v_b_8')
// (2, 30, 'sp4_r_v_b_41')
// (2, 31, 'sp4_r_v_b_28')
// (2, 32, 'neigh_op_tnr_2')
// (2, 32, 'neigh_op_tnr_6')
// (2, 32, 'sp4_r_v_b_17')
// (3, 15, 'sp12_h_r_0')
// (3, 15, 'sp12_v_t_23')
// (3, 16, 'sp12_v_b_23')
// (3, 17, 'sp12_v_b_20')
// (3, 17, 'sp4_h_r_3')
// (3, 17, 'sp4_v_t_47')
// (3, 18, 'sp12_v_b_19')
// (3, 18, 'sp4_v_b_47')
// (3, 19, 'sp12_v_b_16')
// (3, 19, 'sp4_h_r_9')
// (3, 19, 'sp4_v_b_34')
// (3, 19, 'sp4_v_t_41')
// (3, 20, 'sp12_v_b_15')
// (3, 20, 'sp4_v_b_23')
// (3, 20, 'sp4_v_b_41')
// (3, 21, 'sp12_v_b_12')
// (3, 21, 'sp4_h_r_10')
// (3, 21, 'sp4_v_b_10')
// (3, 21, 'sp4_v_b_28')
// (3, 21, 'sp4_v_t_47')
// (3, 22, 'sp12_v_b_11')
// (3, 22, 'sp4_v_b_17')
// (3, 22, 'sp4_v_b_47')
// (3, 23, 'sp12_h_r_0')
// (3, 23, 'sp12_v_b_8')
// (3, 23, 'sp12_v_t_23')
// (3, 23, 'sp4_v_b_34')
// (3, 23, 'sp4_v_b_4')
// (3, 23, 'sp4_v_t_45')
// (3, 24, 'sp12_v_b_23')
// (3, 24, 'sp12_v_b_7')
// (3, 24, 'sp4_v_b_23')
// (3, 24, 'sp4_v_b_45')
// (3, 25, 'sp12_v_b_20')
// (3, 25, 'sp12_v_b_4')
// (3, 25, 'sp4_v_b_10')
// (3, 25, 'sp4_v_b_32')
// (3, 26, 'sp12_v_b_19')
// (3, 26, 'sp12_v_b_3')
// (3, 26, 'sp4_v_b_21')
// (3, 27, 'sp12_h_r_0')
// (3, 27, 'sp12_v_b_0')
// (3, 27, 'sp12_v_b_16')
// (3, 27, 'sp12_v_t_23')
// (3, 27, 'sp4_v_b_8')
// (3, 28, 'sp12_v_b_15')
// (3, 28, 'sp12_v_b_23')
// (3, 29, 'sp12_v_b_12')
// (3, 29, 'sp12_v_b_20')
// (3, 29, 'sp4_h_r_4')
// (3, 29, 'sp4_v_t_41')
// (3, 30, 'sp12_v_b_11')
// (3, 30, 'sp12_v_b_19')
// (3, 30, 'sp4_v_b_41')
// (3, 31, 'sp12_v_b_16')
// (3, 31, 'sp12_v_b_8')
// (3, 31, 'sp4_v_b_28')
// (3, 32, 'neigh_op_top_2')
// (3, 32, 'neigh_op_top_6')
// (3, 32, 'sp12_v_b_15')
// (3, 32, 'sp12_v_b_7')
// (3, 32, 'sp4_v_b_17')
// (3, 33, 'io_1/D_IN_0')
// (3, 33, 'io_1/PAD')
// (3, 33, 'span12_vert_12')
// (3, 33, 'span12_vert_4')
// (3, 33, 'span4_vert_4')
// (4, 15, 'sp12_h_r_3')
// (4, 17, 'sp4_h_r_14')
// (4, 19, 'sp4_h_r_20')
// (4, 21, 'sp4_h_r_23')
// (4, 23, 'sp12_h_r_3')
// (4, 27, 'sp12_h_r_3')
// (4, 29, 'sp4_h_r_17')
// (4, 32, 'neigh_op_tnl_2')
// (4, 32, 'neigh_op_tnl_6')
// (5, 15, 'sp12_h_r_4')
// (5, 17, 'sp4_h_r_27')
// (5, 19, 'sp4_h_r_33')
// (5, 21, 'sp4_h_r_34')
// (5, 23, 'sp12_h_r_4')
// (5, 27, 'sp12_h_r_4')
// (5, 29, 'sp4_h_r_28')
// (6, 15, 'sp12_h_r_7')
// (6, 17, 'sp4_h_r_38')
// (6, 19, 'sp4_h_r_44')
// (6, 21, 'sp4_h_r_47')
// (6, 23, 'sp12_h_r_7')
// (6, 26, 'sp4_r_v_b_41')
// (6, 27, 'sp12_h_r_7')
// (6, 27, 'sp4_r_v_b_28')
// (6, 28, 'sp4_r_v_b_17')
// (6, 29, 'sp4_h_r_41')
// (6, 29, 'sp4_r_v_b_4')
// (7, 15, 'sp12_h_r_8')
// (7, 17, 'sp4_h_l_38')
// (7, 17, 'sp4_h_r_11')
// (7, 19, 'sp4_h_l_44')
// (7, 19, 'sp4_h_r_5')
// (7, 21, 'sp4_h_l_47')
// (7, 21, 'sp4_h_r_10')
// (7, 23, 'sp12_h_r_8')
// (7, 25, 'sp4_h_r_9')
// (7, 25, 'sp4_v_t_41')
// (7, 26, 'sp4_v_b_41')
// (7, 27, 'sp12_h_r_8')
// (7, 27, 'sp4_v_b_28')
// (7, 28, 'sp4_v_b_17')
// (7, 29, 'sp4_h_l_41')
// (7, 29, 'sp4_h_r_4')
// (7, 29, 'sp4_h_r_7')
// (7, 29, 'sp4_v_b_4')
// (8, 15, 'local_g0_3')
// (8, 15, 'ram/RADDR_0')
// (8, 15, 'sp12_h_r_11')
// (8, 17, 'local_g1_6')
// (8, 17, 'ram/RADDR_0')
// (8, 17, 'sp4_h_r_22')
// (8, 19, 'local_g1_0')
// (8, 19, 'ram/RADDR_0')
// (8, 19, 'sp4_h_r_16')
// (8, 21, 'local_g0_7')
// (8, 21, 'ram/RADDR_0')
// (8, 21, 'sp4_h_r_23')
// (8, 23, 'local_g0_7')
// (8, 23, 'ram/RADDR_0')
// (8, 23, 'sp12_h_r_11')
// (8, 23, 'sp4_h_r_7')
// (8, 25, 'local_g1_4')
// (8, 25, 'ram/RADDR_0')
// (8, 25, 'sp4_h_r_20')
// (8, 27, 'local_g0_7')
// (8, 27, 'ram/RADDR_0')
// (8, 27, 'sp12_h_r_11')
// (8, 27, 'sp4_h_r_7')
// (8, 29, 'local_g1_2')
// (8, 29, 'ram/RADDR_0')
// (8, 29, 'sp4_h_r_17')
// (8, 29, 'sp4_h_r_18')
// (9, 15, 'sp12_h_r_12')
// (9, 17, 'sp4_h_r_35')
// (9, 19, 'sp4_h_r_29')
// (9, 21, 'sp4_h_r_34')
// (9, 23, 'sp12_h_r_12')
// (9, 23, 'sp4_h_r_18')
// (9, 25, 'sp4_h_r_33')
// (9, 27, 'sp12_h_r_12')
// (9, 27, 'sp4_h_r_18')
// (9, 29, 'sp4_h_r_28')
// (9, 29, 'sp4_h_r_31')
// (10, 15, 'sp12_h_r_15')
// (10, 17, 'sp4_h_r_46')
// (10, 19, 'sp4_h_r_40')
// (10, 21, 'sp4_h_r_47')
// (10, 23, 'sp12_h_r_15')
// (10, 23, 'sp4_h_r_31')
// (10, 25, 'sp4_h_r_44')
// (10, 27, 'sp12_h_r_15')
// (10, 27, 'sp4_h_r_31')
// (10, 29, 'sp4_h_r_41')
// (10, 29, 'sp4_h_r_42')
// (11, 15, 'sp12_h_r_16')
// (11, 17, 'sp4_h_l_46')
// (11, 19, 'sp4_h_l_40')
// (11, 21, 'sp4_h_l_47')
// (11, 23, 'sp12_h_r_16')
// (11, 23, 'sp4_h_r_42')
// (11, 25, 'sp4_h_l_44')
// (11, 27, 'sp12_h_r_16')
// (11, 27, 'sp4_h_r_42')
// (11, 29, 'sp4_h_l_41')
// (11, 29, 'sp4_h_l_42')
// (11, 29, 'sp4_h_r_7')
// (12, 15, 'sp12_h_r_19')
// (12, 23, 'sp12_h_r_19')
// (12, 23, 'sp4_h_l_42')
// (12, 27, 'sp12_h_r_19')
// (12, 27, 'sp4_h_l_42')
// (12, 29, 'sp4_h_r_18')
// (13, 15, 'sp12_h_r_20')
// (13, 23, 'sp12_h_r_20')
// (13, 27, 'sp12_h_r_20')
// (13, 29, 'sp4_h_r_31')
// (14, 15, 'sp12_h_r_23')
// (14, 23, 'sp12_h_r_23')
// (14, 27, 'sp12_h_r_23')
// (14, 29, 'sp4_h_r_42')
// (15, 15, 'sp12_h_l_23')
// (15, 23, 'sp12_h_l_23')
// (15, 23, 'sp12_h_r_0')
// (15, 27, 'sp12_h_l_23')
// (15, 27, 'sp12_h_r_0')
// (15, 29, 'sp4_h_l_42')
// (15, 29, 'sp4_h_r_10')
// (16, 23, 'sp12_h_r_3')
// (16, 27, 'sp12_h_r_3')
// (16, 29, 'sp4_h_r_23')
// (17, 23, 'sp12_h_r_4')
// (17, 27, 'sp12_h_r_4')
// (17, 29, 'sp4_h_r_34')
// (18, 23, 'sp12_h_r_7')
// (18, 23, 'sp4_h_r_5')
// (18, 27, 'sp12_h_r_7')
// (18, 29, 'sp4_h_r_47')
// (19, 23, 'sp12_h_r_8')
// (19, 23, 'sp4_h_r_16')
// (19, 27, 'sp12_h_r_8')
// (19, 29, 'sp4_h_l_47')
// (19, 29, 'sp4_h_r_10')
// (20, 23, 'sp12_h_r_11')
// (20, 23, 'sp4_h_r_29')
// (20, 23, 'sp4_h_r_7')
// (20, 27, 'sp12_h_r_11')
// (20, 29, 'sp4_h_r_23')
// (21, 16, 'sp4_r_v_b_45')
// (21, 17, 'sp4_r_v_b_32')
// (21, 18, 'sp4_r_v_b_21')
// (21, 19, 'sp4_r_v_b_8')
// (21, 20, 'sp4_r_v_b_40')
// (21, 21, 'sp4_r_v_b_29')
// (21, 22, 'sp4_r_v_b_16')
// (21, 23, 'sp12_h_r_12')
// (21, 23, 'sp4_h_r_18')
// (21, 23, 'sp4_h_r_40')
// (21, 23, 'sp4_r_v_b_5')
// (21, 27, 'sp12_h_r_12')
// (21, 29, 'sp4_h_r_34')
// (22, 15, 'sp4_v_t_45')
// (22, 16, 'sp4_v_b_45')
// (22, 17, 'sp4_v_b_32')
// (22, 18, 'local_g1_5')
// (22, 18, 'lutff_7/in_1')
// (22, 18, 'sp4_v_b_21')
// (22, 19, 'sp4_v_b_8')
// (22, 19, 'sp4_v_t_40')
// (22, 20, 'sp4_v_b_40')
// (22, 21, 'sp4_v_b_29')
// (22, 22, 'sp4_v_b_16')
// (22, 23, 'sp12_h_r_15')
// (22, 23, 'sp4_h_l_40')
// (22, 23, 'sp4_h_r_31')
// (22, 23, 'sp4_h_r_9')
// (22, 23, 'sp4_v_b_5')
// (22, 27, 'sp12_h_r_15')
// (22, 29, 'sp4_h_r_47')
// (23, 16, 'sp4_r_v_b_41')
// (23, 17, 'sp4_r_v_b_28')
// (23, 18, 'sp4_r_v_b_17')
// (23, 19, 'sp4_r_v_b_4')
// (23, 20, 'sp4_r_v_b_36')
// (23, 21, 'local_g1_1')
// (23, 21, 'lutff_6/in_2')
// (23, 21, 'sp4_r_v_b_25')
// (23, 22, 'sp4_r_v_b_12')
// (23, 23, 'sp12_h_r_16')
// (23, 23, 'sp4_h_r_20')
// (23, 23, 'sp4_h_r_42')
// (23, 23, 'sp4_r_v_b_1')
// (23, 27, 'sp12_h_r_16')
// (23, 29, 'sp4_h_l_47')
// (23, 29, 'sp4_h_r_1')
// (24, 15, 'sp4_h_r_4')
// (24, 15, 'sp4_v_t_41')
// (24, 16, 'sp4_v_b_41')
// (24, 17, 'sp4_v_b_28')
// (24, 18, 'sp4_v_b_17')
// (24, 19, 'sp4_h_r_1')
// (24, 19, 'sp4_v_b_4')
// (24, 19, 'sp4_v_t_36')
// (24, 20, 'sp4_v_b_36')
// (24, 21, 'sp4_v_b_25')
// (24, 22, 'sp4_v_b_12')
// (24, 23, 'sp12_h_r_19')
// (24, 23, 'sp4_h_l_42')
// (24, 23, 'sp4_h_r_33')
// (24, 23, 'sp4_v_b_1')
// (24, 27, 'sp12_h_r_19')
// (24, 29, 'sp4_h_r_12')
// (25, 15, 'local_g0_1')
// (25, 15, 'ram/RADDR_0')
// (25, 15, 'sp4_h_r_17')
// (25, 16, 'sp4_r_v_b_38')
// (25, 17, 'local_g0_3')
// (25, 17, 'ram/RADDR_0')
// (25, 17, 'sp4_r_v_b_27')
// (25, 18, 'sp4_r_v_b_14')
// (25, 19, 'local_g1_4')
// (25, 19, 'ram/RADDR_0')
// (25, 19, 'sp4_h_r_12')
// (25, 19, 'sp4_r_v_b_3')
// (25, 20, 'sp4_r_v_b_38')
// (25, 21, 'local_g0_3')
// (25, 21, 'ram/RADDR_0')
// (25, 21, 'sp4_r_v_b_27')
// (25, 22, 'sp4_r_v_b_14')
// (25, 23, 'local_g1_4')
// (25, 23, 'ram/RADDR_0')
// (25, 23, 'sp12_h_r_20')
// (25, 23, 'sp4_h_r_44')
// (25, 23, 'sp4_r_v_b_3')
// (25, 24, 'sp4_r_v_b_39')
// (25, 25, 'local_g1_2')
// (25, 25, 'ram/RADDR_0')
// (25, 25, 'sp4_r_v_b_26')
// (25, 26, 'sp4_r_v_b_15')
// (25, 27, 'local_g1_4')
// (25, 27, 'ram/RADDR_0')
// (25, 27, 'sp12_h_r_20')
// (25, 27, 'sp4_r_v_b_2')
// (25, 29, 'local_g2_1')
// (25, 29, 'ram/RADDR_0')
// (25, 29, 'sp4_h_r_25')
// (26, 15, 'sp4_h_r_28')
// (26, 15, 'sp4_v_t_38')
// (26, 16, 'sp4_v_b_38')
// (26, 17, 'sp4_v_b_27')
// (26, 18, 'sp4_v_b_14')
// (26, 19, 'sp4_h_r_25')
// (26, 19, 'sp4_v_b_3')
// (26, 19, 'sp4_v_t_38')
// (26, 20, 'sp4_v_b_38')
// (26, 21, 'sp4_v_b_27')
// (26, 22, 'sp4_v_b_14')
// (26, 23, 'sp12_h_r_23')
// (26, 23, 'sp4_h_l_44')
// (26, 23, 'sp4_v_b_3')
// (26, 23, 'sp4_v_t_39')
// (26, 24, 'sp4_v_b_39')
// (26, 25, 'sp4_v_b_26')
// (26, 26, 'sp4_v_b_15')
// (26, 27, 'sp12_h_r_23')
// (26, 27, 'sp4_v_b_2')
// (26, 29, 'sp4_h_r_36')
// (27, 15, 'sp4_h_r_41')
// (27, 19, 'sp4_h_r_36')
// (27, 23, 'sp12_h_l_23')
// (27, 27, 'sp12_h_l_23')
// (27, 29, 'sp4_h_l_36')
// (28, 15, 'sp4_h_l_41')
// (28, 19, 'sp4_h_l_36')

wire io_4_33_0;
// (3, 16, 'sp4_r_v_b_43')
// (3, 17, 'sp4_r_v_b_30')
// (3, 18, 'sp4_r_v_b_19')
// (3, 19, 'sp4_r_v_b_6')
// (3, 20, 'sp4_r_v_b_47')
// (3, 21, 'sp4_r_v_b_34')
// (3, 22, 'sp4_r_v_b_23')
// (3, 23, 'sp4_r_v_b_10')
// (3, 26, 'sp4_r_v_b_46')
// (3, 27, 'sp4_r_v_b_35')
// (3, 28, 'sp4_r_v_b_22')
// (3, 29, 'sp4_r_v_b_11')
// (3, 30, 'sp4_r_v_b_45')
// (3, 31, 'sp4_r_v_b_32')
// (3, 32, 'neigh_op_tnr_0')
// (3, 32, 'neigh_op_tnr_4')
// (3, 32, 'sp4_r_v_b_21')
// (4, 15, 'sp4_h_r_11')
// (4, 15, 'sp4_v_t_43')
// (4, 16, 'sp4_v_b_43')
// (4, 17, 'sp4_v_b_30')
// (4, 18, 'sp4_v_b_19')
// (4, 19, 'sp4_h_r_3')
// (4, 19, 'sp4_v_b_6')
// (4, 19, 'sp4_v_t_47')
// (4, 20, 'sp4_v_b_47')
// (4, 21, 'sp12_h_r_0')
// (4, 21, 'sp12_v_t_23')
// (4, 21, 'sp4_v_b_34')
// (4, 22, 'sp12_v_b_23')
// (4, 22, 'sp4_v_b_23')
// (4, 23, 'sp12_v_b_20')
// (4, 23, 'sp4_v_b_10')
// (4, 24, 'sp12_v_b_19')
// (4, 25, 'sp12_h_r_0')
// (4, 25, 'sp12_v_b_16')
// (4, 25, 'sp12_v_t_23')
// (4, 25, 'sp4_h_r_11')
// (4, 25, 'sp4_v_t_46')
// (4, 26, 'sp12_v_b_15')
// (4, 26, 'sp12_v_b_23')
// (4, 26, 'sp4_v_b_46')
// (4, 27, 'sp12_v_b_12')
// (4, 27, 'sp12_v_b_20')
// (4, 27, 'sp4_v_b_35')
// (4, 28, 'sp12_v_b_11')
// (4, 28, 'sp12_v_b_19')
// (4, 28, 'sp4_v_b_22')
// (4, 29, 'sp12_v_b_16')
// (4, 29, 'sp12_v_b_8')
// (4, 29, 'sp4_h_r_1')
// (4, 29, 'sp4_v_b_11')
// (4, 29, 'sp4_v_t_45')
// (4, 30, 'sp12_v_b_15')
// (4, 30, 'sp12_v_b_7')
// (4, 30, 'sp4_v_b_45')
// (4, 31, 'sp12_v_b_12')
// (4, 31, 'sp12_v_b_4')
// (4, 31, 'sp4_v_b_32')
// (4, 32, 'neigh_op_top_0')
// (4, 32, 'neigh_op_top_4')
// (4, 32, 'sp12_v_b_11')
// (4, 32, 'sp12_v_b_3')
// (4, 32, 'sp4_v_b_21')
// (4, 33, 'io_0/D_IN_0')
// (4, 33, 'io_0/PAD')
// (4, 33, 'span12_vert_0')
// (4, 33, 'span12_vert_8')
// (4, 33, 'span4_vert_8')
// (5, 15, 'sp4_h_r_22')
// (5, 19, 'sp4_h_r_14')
// (5, 21, 'sp12_h_r_3')
// (5, 25, 'sp12_h_r_3')
// (5, 25, 'sp4_h_r_22')
// (5, 29, 'sp4_h_r_12')
// (5, 32, 'neigh_op_tnl_0')
// (5, 32, 'neigh_op_tnl_4')
// (6, 15, 'sp4_h_r_35')
// (6, 19, 'sp4_h_r_27')
// (6, 21, 'sp12_h_r_4')
// (6, 25, 'sp12_h_r_4')
// (6, 25, 'sp4_h_r_35')
// (6, 29, 'sp4_h_r_25')
// (7, 15, 'sp4_h_r_46')
// (7, 16, 'sp4_r_v_b_44')
// (7, 17, 'sp4_r_v_b_33')
// (7, 18, 'sp4_r_v_b_20')
// (7, 19, 'sp4_h_r_38')
// (7, 19, 'sp4_r_v_b_9')
// (7, 21, 'sp12_h_r_7')
// (7, 22, 'sp4_r_v_b_40')
// (7, 23, 'sp4_r_v_b_29')
// (7, 24, 'sp4_r_v_b_16')
// (7, 25, 'sp12_h_r_7')
// (7, 25, 'sp4_h_r_46')
// (7, 25, 'sp4_r_v_b_5')
// (7, 26, 'sp4_r_v_b_36')
// (7, 27, 'sp4_r_v_b_25')
// (7, 28, 'sp4_r_v_b_12')
// (7, 29, 'sp4_h_r_36')
// (7, 29, 'sp4_r_v_b_1')
// (8, 15, 'local_g1_7')
// (8, 15, 'ram/RADDR_1')
// (8, 15, 'sp4_h_l_46')
// (8, 15, 'sp4_h_r_7')
// (8, 15, 'sp4_v_t_44')
// (8, 16, 'sp4_v_b_44')
// (8, 17, 'local_g3_1')
// (8, 17, 'ram/RADDR_1')
// (8, 17, 'sp4_v_b_33')
// (8, 18, 'sp4_v_b_20')
// (8, 19, 'local_g1_3')
// (8, 19, 'ram/RADDR_1')
// (8, 19, 'sp4_h_l_38')
// (8, 19, 'sp4_h_r_11')
// (8, 19, 'sp4_v_b_9')
// (8, 21, 'local_g0_0')
// (8, 21, 'ram/RADDR_1')
// (8, 21, 'sp12_h_r_8')
// (8, 21, 'sp4_v_t_40')
// (8, 22, 'sp4_v_b_40')
// (8, 23, 'local_g3_5')
// (8, 23, 'ram/RADDR_1')
// (8, 23, 'sp4_v_b_29')
// (8, 24, 'sp4_v_b_16')
// (8, 25, 'local_g1_7')
// (8, 25, 'ram/RADDR_1')
// (8, 25, 'sp12_h_r_8')
// (8, 25, 'sp4_h_l_46')
// (8, 25, 'sp4_h_r_7')
// (8, 25, 'sp4_v_b_5')
// (8, 25, 'sp4_v_t_36')
// (8, 26, 'sp4_v_b_36')
// (8, 27, 'local_g3_1')
// (8, 27, 'ram/RADDR_1')
// (8, 27, 'sp4_v_b_25')
// (8, 28, 'sp4_v_b_12')
// (8, 29, 'local_g1_1')
// (8, 29, 'ram/RADDR_1')
// (8, 29, 'sp4_h_l_36')
// (8, 29, 'sp4_h_r_1')
// (8, 29, 'sp4_v_b_1')
// (9, 15, 'sp4_h_r_18')
// (9, 19, 'sp4_h_r_22')
// (9, 21, 'sp12_h_r_11')
// (9, 25, 'sp12_h_r_11')
// (9, 25, 'sp4_h_r_18')
// (9, 29, 'sp4_h_r_12')
// (10, 15, 'sp4_h_r_31')
// (10, 19, 'sp4_h_r_35')
// (10, 21, 'sp12_h_r_12')
// (10, 25, 'sp12_h_r_12')
// (10, 25, 'sp4_h_r_31')
// (10, 29, 'sp4_h_r_25')
// (11, 15, 'sp4_h_r_42')
// (11, 19, 'sp4_h_r_46')
// (11, 21, 'sp12_h_r_15')
// (11, 25, 'sp12_h_r_15')
// (11, 25, 'sp4_h_r_42')
// (11, 29, 'sp4_h_r_36')
// (12, 15, 'sp4_h_l_42')
// (12, 19, 'sp4_h_l_46')
// (12, 21, 'sp12_h_r_16')
// (12, 25, 'sp12_h_r_16')
// (12, 25, 'sp4_h_l_42')
// (12, 29, 'sp4_h_l_36')
// (12, 29, 'sp4_h_r_9')
// (13, 21, 'sp12_h_r_19')
// (13, 21, 'sp4_h_r_11')
// (13, 25, 'sp12_h_r_19')
// (13, 29, 'sp4_h_r_20')
// (14, 21, 'sp12_h_r_20')
// (14, 21, 'sp4_h_r_22')
// (14, 25, 'sp12_h_r_20')
// (14, 29, 'sp4_h_r_33')
// (15, 21, 'sp12_h_r_23')
// (15, 21, 'sp4_h_r_35')
// (15, 25, 'sp12_h_r_23')
// (15, 29, 'sp4_h_r_44')
// (16, 21, 'sp12_h_l_23')
// (16, 21, 'sp12_h_r_0')
// (16, 21, 'sp4_h_r_46')
// (16, 25, 'sp12_h_l_23')
// (16, 25, 'sp12_h_r_0')
// (16, 29, 'sp4_h_l_44')
// (16, 29, 'sp4_h_r_9')
// (17, 21, 'sp12_h_r_3')
// (17, 21, 'sp4_h_l_46')
// (17, 21, 'sp4_h_r_11')
// (17, 25, 'sp12_h_r_3')
// (17, 29, 'sp4_h_r_20')
// (18, 21, 'sp12_h_r_4')
// (18, 21, 'sp4_h_r_22')
// (18, 25, 'sp12_h_r_4')
// (18, 29, 'sp4_h_r_33')
// (19, 21, 'sp12_h_r_7')
// (19, 21, 'sp4_h_r_35')
// (19, 25, 'sp12_h_r_7')
// (19, 29, 'sp4_h_r_44')
// (20, 18, 'sp4_r_v_b_40')
// (20, 19, 'sp4_r_v_b_29')
// (20, 20, 'sp4_r_v_b_16')
// (20, 21, 'sp12_h_r_8')
// (20, 21, 'sp4_h_r_46')
// (20, 21, 'sp4_r_v_b_5')
// (20, 25, 'sp12_h_r_8')
// (20, 29, 'sp4_h_l_44')
// (20, 29, 'sp4_h_r_0')
// (21, 17, 'sp4_h_r_5')
// (21, 17, 'sp4_v_t_40')
// (21, 18, 'local_g3_0')
// (21, 18, 'lutff_3/in_2')
// (21, 18, 'sp4_v_b_40')
// (21, 19, 'sp4_v_b_29')
// (21, 20, 'sp4_v_b_16')
// (21, 21, 'sp12_h_r_11')
// (21, 21, 'sp4_h_l_46')
// (21, 21, 'sp4_h_r_2')
// (21, 21, 'sp4_v_b_5')
// (21, 25, 'sp12_h_r_11')
// (21, 29, 'sp4_h_r_13')
// (22, 17, 'sp4_h_r_16')
// (22, 21, 'sp12_h_r_12')
// (22, 21, 'sp4_h_r_15')
// (22, 25, 'sp12_h_r_12')
// (22, 29, 'sp4_h_r_24')
// (23, 17, 'sp4_h_r_29')
// (23, 21, 'local_g1_7')
// (23, 21, 'lutff_6/in_0')
// (23, 21, 'sp12_h_r_15')
// (23, 21, 'sp4_h_r_26')
// (23, 25, 'sp12_h_r_15')
// (23, 29, 'sp4_h_r_37')
// (24, 15, 'sp4_h_r_10')
// (24, 17, 'sp4_h_r_40')
// (24, 18, 'sp4_r_v_b_45')
// (24, 19, 'sp4_r_v_b_32')
// (24, 20, 'sp4_r_v_b_21')
// (24, 21, 'sp12_h_r_16')
// (24, 21, 'sp4_h_r_39')
// (24, 21, 'sp4_r_v_b_8')
// (24, 22, 'sp4_r_v_b_39')
// (24, 23, 'sp4_r_v_b_26')
// (24, 24, 'sp4_r_v_b_15')
// (24, 25, 'sp12_h_r_16')
// (24, 25, 'sp4_r_v_b_2')
// (24, 26, 'sp4_r_v_b_46')
// (24, 27, 'sp4_r_v_b_35')
// (24, 28, 'sp4_r_v_b_22')
// (24, 29, 'sp4_h_l_37')
// (24, 29, 'sp4_h_r_3')
// (24, 29, 'sp4_r_v_b_11')
// (25, 15, 'local_g1_7')
// (25, 15, 'ram/RADDR_1')
// (25, 15, 'sp4_h_r_23')
// (25, 17, 'local_g0_0')
// (25, 17, 'ram/RADDR_1')
// (25, 17, 'sp4_h_l_40')
// (25, 17, 'sp4_h_r_8')
// (25, 17, 'sp4_v_t_45')
// (25, 18, 'sp4_v_b_45')
// (25, 19, 'local_g2_0')
// (25, 19, 'ram/RADDR_1')
// (25, 19, 'sp4_v_b_32')
// (25, 20, 'sp4_v_b_21')
// (25, 21, 'local_g1_3')
// (25, 21, 'ram/RADDR_1')
// (25, 21, 'sp12_h_r_19')
// (25, 21, 'sp4_h_l_39')
// (25, 21, 'sp4_v_b_8')
// (25, 21, 'sp4_v_t_39')
// (25, 22, 'sp4_v_b_39')
// (25, 23, 'local_g2_2')
// (25, 23, 'ram/RADDR_1')
// (25, 23, 'sp4_v_b_26')
// (25, 24, 'sp4_v_b_15')
// (25, 25, 'local_g1_3')
// (25, 25, 'ram/RADDR_1')
// (25, 25, 'sp12_h_r_19')
// (25, 25, 'sp4_h_r_11')
// (25, 25, 'sp4_v_b_2')
// (25, 25, 'sp4_v_t_46')
// (25, 26, 'sp4_v_b_46')
// (25, 27, 'local_g3_3')
// (25, 27, 'ram/RADDR_1')
// (25, 27, 'sp4_v_b_35')
// (25, 28, 'sp4_v_b_22')
// (25, 29, 'local_g0_6')
// (25, 29, 'ram/RADDR_1')
// (25, 29, 'sp4_h_r_14')
// (25, 29, 'sp4_v_b_11')
// (26, 15, 'sp4_h_r_34')
// (26, 17, 'sp4_h_r_21')
// (26, 21, 'sp12_h_r_20')
// (26, 25, 'sp12_h_r_20')
// (26, 25, 'sp4_h_r_22')
// (26, 29, 'sp4_h_r_27')
// (27, 12, 'sp4_r_v_b_47')
// (27, 13, 'sp4_r_v_b_34')
// (27, 14, 'sp4_r_v_b_23')
// (27, 15, 'sp4_h_r_47')
// (27, 15, 'sp4_r_v_b_10')
// (27, 17, 'sp4_h_r_32')
// (27, 21, 'sp12_h_r_23')
// (27, 25, 'sp12_h_r_23')
// (27, 25, 'sp4_h_r_35')
// (27, 29, 'sp4_h_r_38')
// (28, 11, 'sp4_v_t_47')
// (28, 12, 'sp4_v_b_47')
// (28, 13, 'sp12_v_t_23')
// (28, 13, 'sp4_v_b_34')
// (28, 14, 'sp12_v_b_23')
// (28, 14, 'sp4_v_b_23')
// (28, 15, 'sp12_v_b_20')
// (28, 15, 'sp4_h_l_47')
// (28, 15, 'sp4_v_b_10')
// (28, 16, 'sp12_v_b_19')
// (28, 17, 'sp12_v_b_16')
// (28, 17, 'sp4_h_r_45')
// (28, 18, 'sp12_v_b_15')
// (28, 19, 'sp12_v_b_12')
// (28, 20, 'sp12_v_b_11')
// (28, 21, 'sp12_h_l_23')
// (28, 21, 'sp12_v_b_8')
// (28, 22, 'sp12_v_b_7')
// (28, 23, 'sp12_v_b_4')
// (28, 24, 'sp12_v_b_3')
// (28, 25, 'sp12_h_l_23')
// (28, 25, 'sp12_v_b_0')
// (28, 25, 'sp4_h_r_46')
// (28, 29, 'sp4_h_l_38')
// (29, 17, 'sp4_h_l_45')
// (29, 25, 'sp4_h_l_46')

wire n25;
// (3, 17, 'sp12_h_r_1')
// (4, 17, 'sp12_h_r_2')
// (5, 17, 'sp12_h_r_5')
// (6, 17, 'sp12_h_r_6')
// (6, 18, 'sp4_r_v_b_41')
// (6, 19, 'sp4_r_v_b_28')
// (6, 20, 'sp4_r_v_b_17')
// (6, 21, 'sp4_r_v_b_4')
// (7, 17, 'sp12_h_r_9')
// (7, 17, 'sp4_h_r_4')
// (7, 17, 'sp4_v_t_41')
// (7, 18, 'sp4_v_b_41')
// (7, 19, 'sp4_v_b_28')
// (7, 20, 'sp4_v_b_17')
// (7, 21, 'local_g1_4')
// (7, 21, 'lutff_1/in_2')
// (7, 21, 'sp4_v_b_4')
// (8, 17, 'sp12_h_r_10')
// (8, 17, 'sp4_h_r_17')
// (9, 17, 'sp12_h_r_13')
// (9, 17, 'sp4_h_r_28')
// (10, 17, 'sp12_h_r_14')
// (10, 17, 'sp4_h_r_41')
// (11, 17, 'sp12_h_r_17')
// (11, 17, 'sp4_h_l_41')
// (12, 17, 'sp12_h_r_18')
// (13, 17, 'sp12_h_r_21')
// (14, 17, 'sp12_h_r_22')
// (15, 17, 'sp12_h_l_22')
// (15, 17, 'sp12_h_r_1')
// (16, 17, 'sp12_h_r_2')
// (17, 17, 'sp12_h_r_5')
// (18, 17, 'sp12_h_r_6')
// (19, 17, 'sp12_h_r_9')
// (20, 17, 'sp12_h_r_10')
// (21, 17, 'sp12_h_r_13')
// (22, 17, 'sp12_h_r_14')
// (23, 16, 'neigh_op_tnr_5')
// (23, 17, 'neigh_op_rgt_5')
// (23, 17, 'sp12_h_r_17')
// (23, 18, 'neigh_op_bnr_5')
// (24, 16, 'neigh_op_top_5')
// (24, 17, 'lutff_5/out')
// (24, 17, 'sp12_h_r_18')
// (24, 18, 'neigh_op_bot_5')
// (25, 16, 'neigh_op_tnl_5')
// (25, 17, 'neigh_op_lft_5')
// (25, 17, 'sp12_h_r_21')
// (25, 18, 'neigh_op_bnl_5')
// (26, 17, 'sp12_h_r_22')
// (27, 17, 'sp12_h_l_22')

wire io_33_30_1;
// (5, 18, 'sp4_h_r_1')
// (5, 30, 'sp4_h_r_9')
// (6, 18, 'sp4_h_r_12')
// (6, 30, 'sp4_h_r_20')
// (7, 18, 'sp4_h_r_25')
// (7, 30, 'sp4_h_r_33')
// (8, 15, 'local_g3_2')
// (8, 15, 'ram/RADDR_6')
// (8, 15, 'sp4_r_v_b_42')
// (8, 16, 'sp4_r_v_b_31')
// (8, 17, 'local_g3_2')
// (8, 17, 'ram/RADDR_6')
// (8, 17, 'sp4_r_v_b_18')
// (8, 18, 'sp4_h_r_36')
// (8, 18, 'sp4_r_v_b_7')
// (8, 19, 'local_g3_2')
// (8, 19, 'ram/RADDR_6')
// (8, 19, 'sp4_r_v_b_42')
// (8, 20, 'sp4_r_v_b_31')
// (8, 21, 'local_g3_2')
// (8, 21, 'ram/RADDR_6')
// (8, 21, 'sp4_r_v_b_18')
// (8, 22, 'sp4_r_v_b_7')
// (8, 23, 'local_g2_7')
// (8, 23, 'ram/RADDR_6')
// (8, 23, 'sp4_r_v_b_39')
// (8, 24, 'sp4_r_v_b_26')
// (8, 25, 'local_g2_7')
// (8, 25, 'ram/RADDR_6')
// (8, 25, 'sp4_r_v_b_15')
// (8, 26, 'sp4_r_v_b_2')
// (8, 27, 'local_g3_4')
// (8, 27, 'ram/RADDR_6')
// (8, 27, 'sp4_r_v_b_43')
// (8, 27, 'sp4_r_v_b_44')
// (8, 28, 'sp4_r_v_b_30')
// (8, 28, 'sp4_r_v_b_33')
// (8, 29, 'local_g3_4')
// (8, 29, 'ram/RADDR_6')
// (8, 29, 'sp4_r_v_b_19')
// (8, 29, 'sp4_r_v_b_20')
// (8, 30, 'sp4_h_r_44')
// (8, 30, 'sp4_r_v_b_6')
// (8, 30, 'sp4_r_v_b_9')
// (9, 14, 'sp4_v_t_42')
// (9, 15, 'sp4_v_b_42')
// (9, 16, 'sp4_v_b_31')
// (9, 17, 'sp4_v_b_18')
// (9, 18, 'sp4_h_l_36')
// (9, 18, 'sp4_h_r_1')
// (9, 18, 'sp4_v_b_7')
// (9, 18, 'sp4_v_t_42')
// (9, 19, 'sp4_v_b_42')
// (9, 20, 'sp4_v_b_31')
// (9, 21, 'sp4_v_b_18')
// (9, 22, 'sp4_v_b_7')
// (9, 22, 'sp4_v_t_39')
// (9, 23, 'sp4_v_b_39')
// (9, 24, 'sp4_v_b_26')
// (9, 25, 'sp4_v_b_15')
// (9, 26, 'sp4_v_b_2')
// (9, 26, 'sp4_v_t_43')
// (9, 26, 'sp4_v_t_44')
// (9, 27, 'sp4_v_b_43')
// (9, 27, 'sp4_v_b_44')
// (9, 28, 'sp4_v_b_30')
// (9, 28, 'sp4_v_b_33')
// (9, 29, 'sp4_v_b_19')
// (9, 29, 'sp4_v_b_20')
// (9, 30, 'sp4_h_l_44')
// (9, 30, 'sp4_h_r_1')
// (9, 30, 'sp4_v_b_6')
// (9, 30, 'sp4_v_b_9')
// (10, 18, 'sp12_h_r_0')
// (10, 18, 'sp4_h_r_12')
// (10, 30, 'sp12_h_r_0')
// (10, 30, 'sp4_h_r_12')
// (11, 18, 'sp12_h_r_3')
// (11, 18, 'sp4_h_r_25')
// (11, 30, 'sp12_h_r_3')
// (11, 30, 'sp4_h_r_25')
// (12, 18, 'sp12_h_r_4')
// (12, 18, 'sp4_h_r_36')
// (12, 30, 'sp12_h_r_4')
// (12, 30, 'sp4_h_r_36')
// (13, 18, 'sp12_h_r_7')
// (13, 18, 'sp4_h_l_36')
// (13, 30, 'sp12_h_r_7')
// (13, 30, 'sp4_h_l_36')
// (14, 18, 'sp12_h_r_8')
// (14, 30, 'sp12_h_r_8')
// (15, 18, 'sp12_h_r_11')
// (15, 30, 'sp12_h_r_11')
// (16, 18, 'sp12_h_r_12')
// (16, 30, 'sp12_h_r_12')
// (17, 18, 'sp12_h_r_15')
// (17, 30, 'sp12_h_r_15')
// (18, 18, 'sp12_h_r_16')
// (18, 30, 'sp12_h_r_16')
// (19, 18, 'sp12_h_r_19')
// (19, 30, 'sp12_h_r_19')
// (20, 18, 'sp12_h_r_20')
// (20, 30, 'sp12_h_r_20')
// (21, 17, 'sp4_r_v_b_47')
// (21, 18, 'sp12_h_r_23')
// (21, 18, 'sp4_r_v_b_34')
// (21, 19, 'sp4_r_v_b_23')
// (21, 20, 'sp4_r_v_b_10')
// (21, 30, 'sp12_h_r_23')
// (22, 16, 'sp4_h_r_3')
// (22, 16, 'sp4_v_t_47')
// (22, 17, 'sp4_v_b_47')
// (22, 18, 'local_g1_0')
// (22, 18, 'lutff_5/in_0')
// (22, 18, 'sp12_h_l_23')
// (22, 18, 'sp12_h_r_0')
// (22, 18, 'sp12_v_t_23')
// (22, 18, 'sp4_v_b_34')
// (22, 19, 'sp12_v_b_23')
// (22, 19, 'sp4_v_b_23')
// (22, 20, 'sp12_v_b_20')
// (22, 20, 'sp4_v_b_10')
// (22, 21, 'sp12_v_b_19')
// (22, 22, 'local_g3_0')
// (22, 22, 'lutff_6/in_3')
// (22, 22, 'sp12_v_b_16')
// (22, 23, 'sp12_v_b_15')
// (22, 24, 'sp12_v_b_12')
// (22, 25, 'sp12_v_b_11')
// (22, 26, 'sp12_v_b_8')
// (22, 27, 'sp12_v_b_7')
// (22, 28, 'sp12_v_b_4')
// (22, 29, 'sp12_v_b_3')
// (22, 30, 'sp12_h_l_23')
// (22, 30, 'sp12_h_r_0')
// (22, 30, 'sp12_v_b_0')
// (23, 16, 'sp4_h_r_14')
// (23, 18, 'sp12_h_r_3')
// (23, 30, 'sp12_h_r_3')
// (24, 16, 'sp4_h_r_27')
// (24, 18, 'sp12_h_r_4')
// (24, 19, 'sp4_r_v_b_36')
// (24, 20, 'sp4_r_v_b_25')
// (24, 21, 'sp4_r_v_b_12')
// (24, 22, 'sp4_r_v_b_1')
// (24, 23, 'sp4_r_v_b_37')
// (24, 24, 'sp4_r_v_b_24')
// (24, 25, 'sp4_r_v_b_13')
// (24, 26, 'sp4_r_v_b_0')
// (24, 27, 'sp4_r_v_b_43')
// (24, 28, 'sp4_r_v_b_30')
// (24, 29, 'sp4_r_v_b_19')
// (24, 30, 'sp12_h_r_4')
// (24, 30, 'sp4_r_v_b_6')
// (25, 13, 'sp4_r_v_b_44')
// (25, 14, 'sp4_r_v_b_33')
// (25, 15, 'local_g3_4')
// (25, 15, 'ram/RADDR_6')
// (25, 15, 'sp4_r_v_b_20')
// (25, 15, 'sp4_r_v_b_46')
// (25, 16, 'sp4_h_r_38')
// (25, 16, 'sp4_r_v_b_35')
// (25, 16, 'sp4_r_v_b_9')
// (25, 17, 'local_g3_6')
// (25, 17, 'ram/RADDR_6')
// (25, 17, 'sp4_r_v_b_22')
// (25, 18, 'sp12_h_r_7')
// (25, 18, 'sp4_r_v_b_11')
// (25, 18, 'sp4_v_t_36')
// (25, 19, 'sp4_r_v_b_45')
// (25, 19, 'sp4_v_b_36')
// (25, 20, 'sp4_r_v_b_32')
// (25, 20, 'sp4_v_b_25')
// (25, 21, 'local_g1_4')
// (25, 21, 'ram/RADDR_6')
// (25, 21, 'sp4_r_v_b_21')
// (25, 21, 'sp4_v_b_12')
// (25, 22, 'sp4_h_r_1')
// (25, 22, 'sp4_r_v_b_8')
// (25, 22, 'sp4_v_b_1')
// (25, 22, 'sp4_v_t_37')
// (25, 23, 'local_g2_5')
// (25, 23, 'ram/RADDR_6')
// (25, 23, 'sp4_v_b_37')
// (25, 24, 'sp4_v_b_24')
// (25, 25, 'local_g0_5')
// (25, 25, 'ram/RADDR_6')
// (25, 25, 'sp4_v_b_13')
// (25, 26, 'sp4_h_r_7')
// (25, 26, 'sp4_v_b_0')
// (25, 26, 'sp4_v_t_43')
// (25, 27, 'local_g2_3')
// (25, 27, 'ram/RADDR_6')
// (25, 27, 'sp4_v_b_43')
// (25, 28, 'sp4_v_b_30')
// (25, 29, 'local_g0_3')
// (25, 29, 'ram/RADDR_6')
// (25, 29, 'sp4_v_b_19')
// (25, 30, 'sp12_h_r_7')
// (25, 30, 'sp4_h_r_1')
// (25, 30, 'sp4_v_b_6')
// (26, 12, 'sp4_v_t_44')
// (26, 13, 'sp4_v_b_44')
// (26, 14, 'sp4_v_b_33')
// (26, 14, 'sp4_v_t_46')
// (26, 15, 'sp4_v_b_20')
// (26, 15, 'sp4_v_b_46')
// (26, 16, 'sp4_h_l_38')
// (26, 16, 'sp4_v_b_35')
// (26, 16, 'sp4_v_b_9')
// (26, 17, 'sp4_v_b_22')
// (26, 18, 'sp12_h_r_8')
// (26, 18, 'sp12_v_t_23')
// (26, 18, 'sp4_v_b_11')
// (26, 18, 'sp4_v_t_45')
// (26, 19, 'local_g3_7')
// (26, 19, 'lutff_7/in_3')
// (26, 19, 'sp12_v_b_23')
// (26, 19, 'sp4_v_b_45')
// (26, 20, 'sp12_v_b_20')
// (26, 20, 'sp4_v_b_32')
// (26, 21, 'sp12_v_b_19')
// (26, 21, 'sp4_v_b_21')
// (26, 22, 'sp12_v_b_16')
// (26, 22, 'sp4_h_r_12')
// (26, 22, 'sp4_v_b_8')
// (26, 23, 'sp12_v_b_15')
// (26, 24, 'sp12_v_b_12')
// (26, 25, 'sp12_v_b_11')
// (26, 26, 'sp12_v_b_8')
// (26, 26, 'sp4_h_r_18')
// (26, 27, 'sp12_v_b_7')
// (26, 28, 'sp12_v_b_4')
// (26, 29, 'sp12_v_b_3')
// (26, 30, 'sp12_h_r_0')
// (26, 30, 'sp12_h_r_8')
// (26, 30, 'sp12_v_b_0')
// (26, 30, 'sp4_h_r_12')
// (27, 18, 'sp12_h_r_11')
// (27, 22, 'sp4_h_r_25')
// (27, 26, 'sp4_h_r_31')
// (27, 30, 'sp12_h_r_11')
// (27, 30, 'sp12_h_r_3')
// (27, 30, 'sp4_h_r_25')
// (28, 18, 'sp12_h_r_12')
// (28, 22, 'sp4_h_r_36')
// (28, 23, 'sp4_r_v_b_36')
// (28, 24, 'sp4_r_v_b_25')
// (28, 25, 'sp4_r_v_b_12')
// (28, 26, 'sp4_h_r_42')
// (28, 26, 'sp4_r_v_b_1')
// (28, 27, 'sp4_r_v_b_36')
// (28, 28, 'sp4_r_v_b_25')
// (28, 29, 'sp4_r_v_b_12')
// (28, 30, 'sp12_h_r_12')
// (28, 30, 'sp12_h_r_4')
// (28, 30, 'sp4_h_r_36')
// (28, 30, 'sp4_r_v_b_1')
// (29, 18, 'sp12_h_r_15')
// (29, 22, 'sp4_h_l_36')
// (29, 22, 'sp4_v_t_36')
// (29, 23, 'sp4_v_b_36')
// (29, 24, 'sp4_v_b_25')
// (29, 25, 'sp4_v_b_12')
// (29, 26, 'sp4_h_l_42')
// (29, 26, 'sp4_v_b_1')
// (29, 26, 'sp4_v_t_36')
// (29, 27, 'sp4_v_b_36')
// (29, 28, 'sp4_v_b_25')
// (29, 29, 'sp4_v_b_12')
// (29, 30, 'sp12_h_r_15')
// (29, 30, 'sp12_h_r_7')
// (29, 30, 'sp4_h_l_36')
// (29, 30, 'sp4_h_r_1')
// (29, 30, 'sp4_v_b_1')
// (30, 18, 'sp12_h_r_16')
// (30, 30, 'sp12_h_r_16')
// (30, 30, 'sp12_h_r_8')
// (30, 30, 'sp4_h_r_12')
// (31, 18, 'sp12_h_r_19')
// (31, 30, 'sp12_h_r_11')
// (31, 30, 'sp12_h_r_19')
// (31, 30, 'sp4_h_r_25')
// (32, 18, 'sp12_h_r_20')
// (32, 29, 'neigh_op_tnr_2')
// (32, 29, 'neigh_op_tnr_6')
// (32, 30, 'neigh_op_rgt_2')
// (32, 30, 'neigh_op_rgt_6')
// (32, 30, 'sp12_h_r_12')
// (32, 30, 'sp12_h_r_20')
// (32, 30, 'sp4_h_r_36')
// (32, 31, 'neigh_op_bnr_2')
// (32, 31, 'neigh_op_bnr_6')
// (33, 18, 'span12_horz_20')
// (33, 30, 'io_1/D_IN_0')
// (33, 30, 'io_1/PAD')
// (33, 30, 'span12_horz_12')
// (33, 30, 'span12_horz_20')
// (33, 30, 'span4_horz_36')

reg n27 = 0;
// (5, 19, 'neigh_op_tnr_1')
// (5, 20, 'neigh_op_rgt_1')
// (5, 21, 'neigh_op_bnr_1')
// (6, 19, 'neigh_op_top_1')
// (6, 19, 'sp4_r_v_b_46')
// (6, 20, 'local_g0_1')
// (6, 20, 'lutff_1/in_0')
// (6, 20, 'lutff_1/out')
// (6, 20, 'sp4_r_v_b_35')
// (6, 21, 'local_g0_1')
// (6, 21, 'lutff_2/in_1')
// (6, 21, 'neigh_op_bot_1')
// (6, 21, 'sp4_r_v_b_22')
// (6, 22, 'sp4_r_v_b_11')
// (7, 18, 'sp4_v_t_46')
// (7, 19, 'neigh_op_tnl_1')
// (7, 19, 'sp4_v_b_46')
// (7, 20, 'local_g1_1')
// (7, 20, 'lutff_0/in_2')
// (7, 20, 'neigh_op_lft_1')
// (7, 20, 'sp4_v_b_35')
// (7, 21, 'neigh_op_bnl_1')
// (7, 21, 'sp4_v_b_22')
// (7, 22, 'local_g1_3')
// (7, 22, 'lutff_1/in_1')
// (7, 22, 'sp4_v_b_11')

wire n28;
// (5, 19, 'sp12_h_r_0')
// (6, 19, 'sp12_h_r_3')
// (7, 19, 'sp12_h_r_4')
// (8, 19, 'sp12_h_r_7')
// (9, 19, 'local_g0_0')
// (9, 19, 'lutff_0/in_0')
// (9, 19, 'sp12_h_r_8')
// (10, 19, 'sp12_h_r_11')
// (11, 19, 'sp12_h_r_12')
// (12, 19, 'sp12_h_r_15')
// (13, 19, 'sp12_h_r_16')
// (14, 19, 'sp12_h_r_19')
// (15, 19, 'sp12_h_r_20')
// (16, 19, 'sp12_h_r_23')
// (17, 19, 'sp12_h_l_23')
// (17, 19, 'sp12_h_r_0')
// (18, 19, 'sp12_h_r_3')
// (19, 19, 'sp12_h_r_4')
// (20, 19, 'sp12_h_r_7')
// (21, 19, 'sp12_h_r_8')
// (22, 19, 'sp12_h_r_11')
// (23, 19, 'sp12_h_r_12')
// (24, 18, 'neigh_op_tnr_4')
// (24, 19, 'neigh_op_rgt_4')
// (24, 19, 'sp12_h_r_15')
// (24, 20, 'neigh_op_bnr_4')
// (25, 18, 'neigh_op_top_4')
// (25, 19, 'ram/RDATA_11')
// (25, 19, 'sp12_h_r_16')
// (25, 20, 'neigh_op_bot_4')
// (26, 18, 'neigh_op_tnl_4')
// (26, 19, 'neigh_op_lft_4')
// (26, 19, 'sp12_h_r_19')
// (26, 20, 'neigh_op_bnl_4')
// (27, 19, 'sp12_h_r_20')
// (28, 19, 'sp12_h_r_23')
// (29, 19, 'sp12_h_l_23')

wire io_30_33_1;
// (5, 19, 'sp4_h_r_11')
// (6, 11, 'sp12_h_r_0')
// (6, 19, 'sp4_h_r_22')
// (6, 23, 'sp12_h_r_0')
// (6, 29, 'sp4_h_r_11')
// (7, 11, 'sp12_h_r_3')
// (7, 19, 'sp4_h_r_35')
// (7, 23, 'sp12_h_r_3')
// (7, 29, 'sp4_h_r_22')
// (8, 11, 'sp12_h_r_4')
// (8, 12, 'sp4_r_v_b_46')
// (8, 13, 'sp4_r_v_b_35')
// (8, 14, 'sp4_r_v_b_22')
// (8, 15, 'local_g2_3')
// (8, 15, 'ram/RADDR_2')
// (8, 15, 'sp4_r_v_b_11')
// (8, 16, 'sp4_r_v_b_36')
// (8, 17, 'local_g0_1')
// (8, 17, 'ram/RADDR_2')
// (8, 17, 'sp4_r_v_b_25')
// (8, 18, 'sp4_r_v_b_12')
// (8, 19, 'local_g3_6')
// (8, 19, 'ram/RADDR_2')
// (8, 19, 'sp4_h_r_46')
// (8, 19, 'sp4_r_v_b_1')
// (8, 20, 'sp4_r_v_b_40')
// (8, 21, 'local_g0_5')
// (8, 21, 'ram/RADDR_2')
// (8, 21, 'sp4_r_v_b_29')
// (8, 22, 'sp4_r_v_b_16')
// (8, 23, 'local_g1_4')
// (8, 23, 'ram/RADDR_2')
// (8, 23, 'sp12_h_r_4')
// (8, 23, 'sp4_r_v_b_5')
// (8, 24, 'sp4_r_v_b_40')
// (8, 24, 'sp4_r_v_b_46')
// (8, 25, 'local_g0_5')
// (8, 25, 'ram/RADDR_2')
// (8, 25, 'sp4_r_v_b_29')
// (8, 25, 'sp4_r_v_b_35')
// (8, 26, 'sp4_r_v_b_16')
// (8, 26, 'sp4_r_v_b_22')
// (8, 27, 'local_g2_3')
// (8, 27, 'ram/RADDR_2')
// (8, 27, 'sp4_r_v_b_11')
// (8, 27, 'sp4_r_v_b_5')
// (8, 29, 'local_g2_3')
// (8, 29, 'ram/RADDR_2')
// (8, 29, 'sp4_h_r_35')
// (9, 11, 'sp12_h_r_7')
// (9, 11, 'sp4_h_r_5')
// (9, 11, 'sp4_v_t_46')
// (9, 12, 'sp4_v_b_46')
// (9, 13, 'sp4_v_b_35')
// (9, 14, 'sp4_v_b_22')
// (9, 15, 'sp4_v_b_11')
// (9, 15, 'sp4_v_t_36')
// (9, 16, 'sp4_v_b_36')
// (9, 17, 'sp4_v_b_25')
// (9, 18, 'sp4_v_b_12')
// (9, 19, 'sp4_h_l_46')
// (9, 19, 'sp4_v_b_1')
// (9, 19, 'sp4_v_t_40')
// (9, 20, 'sp4_v_b_40')
// (9, 21, 'sp4_v_b_29')
// (9, 22, 'sp4_v_b_16')
// (9, 23, 'sp12_h_r_7')
// (9, 23, 'sp4_h_r_5')
// (9, 23, 'sp4_v_b_5')
// (9, 23, 'sp4_v_t_40')
// (9, 23, 'sp4_v_t_46')
// (9, 24, 'sp4_v_b_40')
// (9, 24, 'sp4_v_b_46')
// (9, 25, 'sp4_v_b_29')
// (9, 25, 'sp4_v_b_35')
// (9, 26, 'sp4_v_b_16')
// (9, 26, 'sp4_v_b_22')
// (9, 27, 'sp4_v_b_11')
// (9, 27, 'sp4_v_b_5')
// (9, 29, 'sp4_h_r_46')
// (10, 11, 'sp12_h_r_8')
// (10, 11, 'sp4_h_r_16')
// (10, 23, 'sp12_h_r_8')
// (10, 23, 'sp4_h_r_16')
// (10, 29, 'sp4_h_l_46')
// (10, 29, 'sp4_h_r_3')
// (11, 11, 'sp12_h_r_11')
// (11, 11, 'sp4_h_r_29')
// (11, 23, 'sp12_h_r_11')
// (11, 23, 'sp4_h_r_29')
// (11, 29, 'sp4_h_r_14')
// (12, 11, 'sp12_h_r_12')
// (12, 11, 'sp4_h_r_40')
// (12, 23, 'sp12_h_r_12')
// (12, 23, 'sp4_h_r_40')
// (12, 29, 'sp4_h_r_27')
// (13, 11, 'sp12_h_r_15')
// (13, 11, 'sp4_h_l_40')
// (13, 23, 'sp12_h_r_15')
// (13, 23, 'sp4_h_l_40')
// (13, 29, 'sp4_h_r_38')
// (14, 11, 'sp12_h_r_16')
// (14, 23, 'sp12_h_r_16')
// (14, 29, 'sp4_h_l_38')
// (14, 29, 'sp4_h_r_0')
// (15, 11, 'sp12_h_r_19')
// (15, 23, 'sp12_h_r_19')
// (15, 29, 'sp4_h_r_13')
// (16, 11, 'sp12_h_r_20')
// (16, 23, 'sp12_h_r_20')
// (16, 29, 'sp4_h_r_24')
// (17, 11, 'sp12_h_r_23')
// (17, 23, 'sp12_h_r_23')
// (17, 29, 'sp4_h_r_37')
// (18, 11, 'sp12_h_l_23')
// (18, 11, 'sp12_v_t_23')
// (18, 12, 'sp12_v_b_23')
// (18, 13, 'sp12_v_b_20')
// (18, 14, 'sp12_v_b_19')
// (18, 15, 'sp12_v_b_16')
// (18, 16, 'sp12_v_b_15')
// (18, 17, 'sp12_v_b_12')
// (18, 18, 'sp12_v_b_11')
// (18, 19, 'sp12_v_b_8')
// (18, 20, 'sp12_v_b_7')
// (18, 21, 'sp12_v_b_4')
// (18, 22, 'sp12_v_b_3')
// (18, 23, 'sp12_h_l_23')
// (18, 23, 'sp12_h_r_0')
// (18, 23, 'sp12_v_b_0')
// (18, 29, 'sp4_h_l_37')
// (18, 29, 'sp4_h_r_0')
// (19, 23, 'sp12_h_r_3')
// (19, 29, 'sp4_h_r_13')
// (20, 23, 'sp12_h_r_4')
// (20, 29, 'sp4_h_r_24')
// (21, 18, 'sp4_r_v_b_36')
// (21, 19, 'sp4_r_v_b_25')
// (21, 20, 'sp4_r_v_b_12')
// (21, 21, 'sp4_r_v_b_1')
// (21, 23, 'sp12_h_r_7')
// (21, 29, 'sp4_h_r_37')
// (22, 17, 'sp4_v_t_36')
// (22, 18, 'local_g3_4')
// (22, 18, 'lutff_0/in_3')
// (22, 18, 'sp4_v_b_36')
// (22, 19, 'sp4_v_b_25')
// (22, 20, 'sp4_v_b_12')
// (22, 21, 'sp4_h_r_1')
// (22, 21, 'sp4_v_b_1')
// (22, 23, 'sp12_h_r_8')
// (22, 29, 'sp4_h_l_37')
// (22, 29, 'sp4_h_r_0')
// (23, 21, 'local_g1_4')
// (23, 21, 'lutff_6/in_1')
// (23, 21, 'sp4_h_r_12')
// (23, 23, 'sp12_h_r_11')
// (23, 29, 'sp4_h_r_13')
// (24, 21, 'sp4_h_r_25')
// (24, 23, 'sp12_h_r_12')
// (24, 29, 'sp4_h_r_24')
// (25, 12, 'sp4_r_v_b_43')
// (25, 13, 'sp4_r_v_b_30')
// (25, 14, 'sp4_r_v_b_19')
// (25, 14, 'sp4_r_v_b_43')
// (25, 15, 'local_g1_6')
// (25, 15, 'ram/RADDR_2')
// (25, 15, 'sp4_r_v_b_30')
// (25, 15, 'sp4_r_v_b_6')
// (25, 16, 'sp4_r_v_b_19')
// (25, 17, 'local_g1_6')
// (25, 17, 'ram/RADDR_2')
// (25, 17, 'sp4_r_v_b_6')
// (25, 18, 'sp4_r_v_b_47')
// (25, 19, 'local_g0_1')
// (25, 19, 'ram/RADDR_2')
// (25, 19, 'sp4_r_v_b_34')
// (25, 20, 'sp4_r_v_b_23')
// (25, 21, 'local_g3_4')
// (25, 21, 'ram/RADDR_2')
// (25, 21, 'sp4_h_r_36')
// (25, 21, 'sp4_r_v_b_10')
// (25, 22, 'sp4_r_v_b_37')
// (25, 23, 'local_g0_7')
// (25, 23, 'ram/RADDR_2')
// (25, 23, 'sp12_h_r_15')
// (25, 23, 'sp4_r_v_b_24')
// (25, 24, 'sp4_r_v_b_13')
// (25, 25, 'local_g1_0')
// (25, 25, 'ram/RADDR_2')
// (25, 25, 'sp4_r_v_b_0')
// (25, 26, 'sp4_r_v_b_41')
// (25, 26, 'sp4_r_v_b_44')
// (25, 27, 'local_g2_1')
// (25, 27, 'ram/RADDR_2')
// (25, 27, 'sp4_r_v_b_28')
// (25, 27, 'sp4_r_v_b_33')
// (25, 28, 'sp4_r_v_b_17')
// (25, 28, 'sp4_r_v_b_20')
// (25, 29, 'local_g1_4')
// (25, 29, 'ram/RADDR_2')
// (25, 29, 'sp4_h_r_37')
// (25, 29, 'sp4_r_v_b_4')
// (25, 29, 'sp4_r_v_b_9')
// (26, 11, 'sp4_v_t_43')
// (26, 12, 'sp4_v_b_43')
// (26, 13, 'sp4_v_b_30')
// (26, 13, 'sp4_v_t_43')
// (26, 14, 'sp4_v_b_19')
// (26, 14, 'sp4_v_b_43')
// (26, 15, 'sp4_h_r_1')
// (26, 15, 'sp4_v_b_30')
// (26, 15, 'sp4_v_b_6')
// (26, 16, 'sp4_v_b_19')
// (26, 17, 'sp4_v_b_6')
// (26, 17, 'sp4_v_t_47')
// (26, 18, 'sp4_v_b_47')
// (26, 19, 'sp4_v_b_34')
// (26, 20, 'sp4_v_b_23')
// (26, 21, 'sp4_h_l_36')
// (26, 21, 'sp4_h_r_10')
// (26, 21, 'sp4_v_b_10')
// (26, 21, 'sp4_v_t_37')
// (26, 22, 'sp4_v_b_37')
// (26, 23, 'sp12_h_r_16')
// (26, 23, 'sp4_v_b_24')
// (26, 24, 'sp4_v_b_13')
// (26, 25, 'sp4_h_r_7')
// (26, 25, 'sp4_v_b_0')
// (26, 25, 'sp4_v_t_41')
// (26, 25, 'sp4_v_t_44')
// (26, 26, 'sp4_v_b_41')
// (26, 26, 'sp4_v_b_44')
// (26, 27, 'sp4_v_b_28')
// (26, 27, 'sp4_v_b_33')
// (26, 28, 'sp4_v_b_17')
// (26, 28, 'sp4_v_b_20')
// (26, 29, 'sp4_h_l_37')
// (26, 29, 'sp4_h_r_4')
// (26, 29, 'sp4_v_b_4')
// (26, 29, 'sp4_v_b_9')
// (27, 15, 'sp4_h_r_12')
// (27, 21, 'sp4_h_r_23')
// (27, 23, 'sp12_h_r_19')
// (27, 25, 'sp4_h_r_18')
// (27, 29, 'sp4_h_r_17')
// (28, 15, 'sp4_h_r_25')
// (28, 21, 'sp4_h_r_34')
// (28, 23, 'sp12_h_r_20')
// (28, 25, 'sp4_h_r_31')
// (28, 29, 'sp4_h_r_28')
// (29, 12, 'sp4_r_v_b_45')
// (29, 13, 'sp4_r_v_b_32')
// (29, 14, 'sp4_r_v_b_21')
// (29, 15, 'sp4_h_r_36')
// (29, 15, 'sp4_r_v_b_8')
// (29, 21, 'sp4_h_r_47')
// (29, 22, 'sp4_r_v_b_47')
// (29, 23, 'sp12_h_r_23')
// (29, 23, 'sp4_r_v_b_34')
// (29, 24, 'sp4_r_v_b_23')
// (29, 25, 'sp4_h_r_42')
// (29, 25, 'sp4_r_v_b_10')
// (29, 26, 'sp4_r_v_b_42')
// (29, 27, 'sp4_r_v_b_31')
// (29, 28, 'sp4_r_v_b_18')
// (29, 29, 'sp4_h_r_41')
// (29, 29, 'sp4_r_v_b_7')
// (29, 30, 'sp4_r_v_b_41')
// (29, 31, 'sp4_r_v_b_28')
// (29, 32, 'neigh_op_tnr_2')
// (29, 32, 'neigh_op_tnr_6')
// (29, 32, 'sp4_r_v_b_17')
// (30, 11, 'sp12_v_t_23')
// (30, 11, 'sp4_v_t_45')
// (30, 12, 'sp12_v_b_23')
// (30, 12, 'sp4_v_b_45')
// (30, 13, 'sp12_v_b_20')
// (30, 13, 'sp4_v_b_32')
// (30, 14, 'sp12_v_b_19')
// (30, 14, 'sp4_v_b_21')
// (30, 15, 'sp12_v_b_16')
// (30, 15, 'sp4_h_l_36')
// (30, 15, 'sp4_v_b_8')
// (30, 16, 'sp12_v_b_15')
// (30, 17, 'sp12_v_b_12')
// (30, 18, 'sp12_v_b_11')
// (30, 19, 'sp12_v_b_8')
// (30, 20, 'sp12_v_b_7')
// (30, 21, 'sp12_v_b_4')
// (30, 21, 'sp4_h_l_47')
// (30, 21, 'sp4_v_t_47')
// (30, 22, 'sp12_v_b_3')
// (30, 22, 'sp4_v_b_47')
// (30, 23, 'sp12_h_l_23')
// (30, 23, 'sp12_v_b_0')
// (30, 23, 'sp12_v_t_23')
// (30, 23, 'sp4_v_b_34')
// (30, 24, 'sp12_v_b_23')
// (30, 24, 'sp4_v_b_23')
// (30, 25, 'sp12_v_b_20')
// (30, 25, 'sp4_h_l_42')
// (30, 25, 'sp4_v_b_10')
// (30, 25, 'sp4_v_t_42')
// (30, 26, 'sp12_v_b_19')
// (30, 26, 'sp4_v_b_42')
// (30, 27, 'sp12_v_b_16')
// (30, 27, 'sp4_v_b_31')
// (30, 28, 'sp12_v_b_15')
// (30, 28, 'sp4_v_b_18')
// (30, 29, 'sp12_v_b_12')
// (30, 29, 'sp4_h_l_41')
// (30, 29, 'sp4_v_b_7')
// (30, 29, 'sp4_v_t_41')
// (30, 30, 'sp12_v_b_11')
// (30, 30, 'sp4_v_b_41')
// (30, 31, 'sp12_v_b_8')
// (30, 31, 'sp4_v_b_28')
// (30, 32, 'neigh_op_top_2')
// (30, 32, 'neigh_op_top_6')
// (30, 32, 'sp12_v_b_7')
// (30, 32, 'sp4_v_b_17')
// (30, 33, 'io_1/D_IN_0')
// (30, 33, 'io_1/PAD')
// (30, 33, 'span12_vert_4')
// (30, 33, 'span4_vert_4')
// (31, 32, 'neigh_op_tnl_2')
// (31, 32, 'neigh_op_tnl_6')

wire n30;
// (5, 19, 'sp4_h_r_6')
// (6, 19, 'sp4_h_r_19')
// (6, 23, 'sp4_h_r_3')
// (7, 19, 'local_g2_6')
// (7, 19, 'local_g3_6')
// (7, 19, 'lutff_2/in_0')
// (7, 19, 'lutff_4/in_1')
// (7, 19, 'sp4_h_r_30')
// (7, 20, 'sp4_r_v_b_41')
// (7, 21, 'local_g0_4')
// (7, 21, 'lutff_2/in_0')
// (7, 21, 'lutff_6/in_2')
// (7, 21, 'sp4_r_v_b_28')
// (7, 22, 'sp4_r_v_b_17')
// (7, 23, 'local_g0_6')
// (7, 23, 'local_g1_6')
// (7, 23, 'lutff_0/in_3')
// (7, 23, 'lutff_6/in_2')
// (7, 23, 'sp4_h_r_14')
// (7, 23, 'sp4_r_v_b_4')
// (7, 24, 'sp4_r_v_b_46')
// (7, 25, 'local_g0_0')
// (7, 25, 'lutff_0/in_2')
// (7, 25, 'sp4_r_v_b_35')
// (7, 26, 'sp4_r_v_b_22')
// (7, 27, 'sp4_r_v_b_11')
// (8, 19, 'sp4_h_r_43')
// (8, 19, 'sp4_v_t_41')
// (8, 20, 'sp4_r_v_b_43')
// (8, 20, 'sp4_v_b_41')
// (8, 21, 'sp4_r_v_b_30')
// (8, 21, 'sp4_v_b_28')
// (8, 22, 'neigh_op_tnr_3')
// (8, 22, 'sp4_r_v_b_19')
// (8, 22, 'sp4_v_b_17')
// (8, 23, 'neigh_op_rgt_3')
// (8, 23, 'sp4_h_r_11')
// (8, 23, 'sp4_h_r_27')
// (8, 23, 'sp4_r_v_b_38')
// (8, 23, 'sp4_r_v_b_6')
// (8, 23, 'sp4_v_b_4')
// (8, 23, 'sp4_v_t_46')
// (8, 24, 'neigh_op_bnr_3')
// (8, 24, 'sp4_r_v_b_27')
// (8, 24, 'sp4_v_b_46')
// (8, 25, 'sp4_r_v_b_14')
// (8, 25, 'sp4_v_b_35')
// (8, 26, 'sp4_r_v_b_3')
// (8, 26, 'sp4_v_b_22')
// (8, 27, 'sp4_v_b_11')
// (9, 19, 'sp4_h_l_43')
// (9, 19, 'sp4_v_t_43')
// (9, 20, 'sp4_v_b_43')
// (9, 21, 'sp4_v_b_30')
// (9, 22, 'neigh_op_top_3')
// (9, 22, 'sp4_v_b_19')
// (9, 22, 'sp4_v_t_38')
// (9, 23, 'lutff_3/out')
// (9, 23, 'sp4_h_r_22')
// (9, 23, 'sp4_h_r_38')
// (9, 23, 'sp4_v_b_38')
// (9, 23, 'sp4_v_b_6')
// (9, 24, 'neigh_op_bot_3')
// (9, 24, 'sp4_v_b_27')
// (9, 25, 'local_g0_6')
// (9, 25, 'lutff_6/in_0')
// (9, 25, 'sp4_v_b_14')
// (9, 26, 'sp4_v_b_3')
// (10, 22, 'neigh_op_tnl_3')
// (10, 23, 'neigh_op_lft_3')
// (10, 23, 'sp4_h_l_38')
// (10, 23, 'sp4_h_r_35')
// (10, 24, 'neigh_op_bnl_3')
// (11, 23, 'sp4_h_r_46')
// (12, 23, 'sp4_h_l_46')

wire n31;
// (5, 20, 'neigh_op_tnr_2')
// (5, 21, 'neigh_op_rgt_2')
// (5, 22, 'neigh_op_bnr_2')
// (6, 20, 'neigh_op_top_2')
// (6, 21, 'local_g0_2')
// (6, 21, 'lutff_2/out')
// (6, 21, 'lutff_global/cen')
// (6, 22, 'neigh_op_bot_2')
// (7, 20, 'neigh_op_tnl_2')
// (7, 21, 'neigh_op_lft_2')
// (7, 22, 'neigh_op_bnl_2')

reg n32 = 0;
// (5, 20, 'neigh_op_tnr_3')
// (5, 21, 'neigh_op_rgt_3')
// (5, 22, 'neigh_op_bnr_3')
// (6, 20, 'neigh_op_top_3')
// (6, 21, 'local_g3_3')
// (6, 21, 'lutff_3/in_1')
// (6, 21, 'lutff_3/out')
// (6, 22, 'neigh_op_bot_3')
// (7, 20, 'local_g3_3')
// (7, 20, 'lutff_1/in_1')
// (7, 20, 'neigh_op_tnl_3')
// (7, 21, 'local_g1_3')
// (7, 21, 'lutff_1/in_3')
// (7, 21, 'neigh_op_lft_3')
// (7, 22, 'neigh_op_bnl_3')

wire n33;
// (5, 22, 'sp4_h_r_1')
// (6, 22, 'sp4_h_r_12')
// (7, 22, 'local_g3_1')
// (7, 22, 'lutff_5/in_3')
// (7, 22, 'sp4_h_r_25')
// (8, 22, 'sp4_h_r_36')
// (8, 23, 'sp4_r_v_b_36')
// (8, 24, 'neigh_op_tnr_6')
// (8, 24, 'sp4_r_v_b_25')
// (8, 25, 'neigh_op_rgt_6')
// (8, 25, 'sp4_r_v_b_12')
// (8, 26, 'neigh_op_bnr_6')
// (8, 26, 'sp4_r_v_b_1')
// (9, 22, 'sp4_h_l_36')
// (9, 22, 'sp4_v_t_36')
// (9, 23, 'sp4_v_b_36')
// (9, 24, 'neigh_op_top_6')
// (9, 24, 'sp4_v_b_25')
// (9, 25, 'lutff_6/out')
// (9, 25, 'sp4_v_b_12')
// (9, 26, 'neigh_op_bot_6')
// (9, 26, 'sp4_v_b_1')
// (10, 24, 'neigh_op_tnl_6')
// (10, 25, 'neigh_op_lft_6')
// (10, 26, 'neigh_op_bnl_6')

wire io_31_33_0;
// (6, 12, 'sp4_r_v_b_43')
// (6, 13, 'sp4_r_v_b_30')
// (6, 14, 'sp4_r_v_b_19')
// (6, 15, 'sp4_r_v_b_6')
// (6, 21, 'sp4_h_r_1')
// (7, 9, 'sp12_v_t_23')
// (7, 10, 'sp12_v_b_23')
// (7, 11, 'sp12_v_b_20')
// (7, 11, 'sp4_v_t_43')
// (7, 12, 'sp12_v_b_19')
// (7, 12, 'sp4_v_b_43')
// (7, 13, 'sp12_v_b_16')
// (7, 13, 'sp4_v_b_30')
// (7, 14, 'sp12_v_b_15')
// (7, 14, 'sp4_v_b_19')
// (7, 15, 'sp12_v_b_12')
// (7, 15, 'sp4_h_r_6')
// (7, 15, 'sp4_v_b_6')
// (7, 16, 'sp12_v_b_11')
// (7, 17, 'sp12_v_b_8')
// (7, 18, 'sp12_v_b_7')
// (7, 18, 'sp4_r_v_b_38')
// (7, 19, 'sp12_v_b_4')
// (7, 19, 'sp4_r_v_b_27')
// (7, 20, 'sp12_v_b_3')
// (7, 20, 'sp4_r_v_b_14')
// (7, 21, 'sp12_h_r_0')
// (7, 21, 'sp12_v_b_0')
// (7, 21, 'sp4_h_r_12')
// (7, 21, 'sp4_r_v_b_3')
// (7, 22, 'sp4_r_v_b_38')
// (7, 22, 'sp4_r_v_b_44')
// (7, 23, 'sp4_r_v_b_27')
// (7, 23, 'sp4_r_v_b_33')
// (7, 24, 'sp4_r_v_b_14')
// (7, 24, 'sp4_r_v_b_20')
// (7, 25, 'sp4_r_v_b_3')
// (7, 25, 'sp4_r_v_b_9')
// (7, 26, 'sp4_r_v_b_43')
// (7, 27, 'sp4_r_v_b_30')
// (7, 28, 'sp4_r_v_b_19')
// (7, 29, 'sp4_r_v_b_6')
// (8, 15, 'local_g1_3')
// (8, 15, 'ram/RADDR_5')
// (8, 15, 'sp4_h_r_19')
// (8, 17, 'local_g1_3')
// (8, 17, 'ram/RADDR_5')
// (8, 17, 'sp4_h_r_3')
// (8, 17, 'sp4_v_t_38')
// (8, 18, 'sp4_v_b_38')
// (8, 19, 'local_g3_3')
// (8, 19, 'ram/RADDR_5')
// (8, 19, 'sp4_v_b_27')
// (8, 20, 'sp4_v_b_14')
// (8, 21, 'local_g3_1')
// (8, 21, 'ram/RADDR_5')
// (8, 21, 'sp12_h_r_3')
// (8, 21, 'sp4_h_r_25')
// (8, 21, 'sp4_h_r_3')
// (8, 21, 'sp4_v_b_3')
// (8, 21, 'sp4_v_t_38')
// (8, 21, 'sp4_v_t_44')
// (8, 22, 'sp4_v_b_38')
// (8, 22, 'sp4_v_b_44')
// (8, 23, 'local_g3_3')
// (8, 23, 'ram/RADDR_5')
// (8, 23, 'sp4_v_b_27')
// (8, 23, 'sp4_v_b_33')
// (8, 24, 'sp4_v_b_14')
// (8, 24, 'sp4_v_b_20')
// (8, 25, 'local_g1_1')
// (8, 25, 'ram/RADDR_5')
// (8, 25, 'sp4_v_b_3')
// (8, 25, 'sp4_v_b_9')
// (8, 25, 'sp4_v_t_43')
// (8, 26, 'sp4_v_b_43')
// (8, 27, 'local_g2_6')
// (8, 27, 'ram/RADDR_5')
// (8, 27, 'sp4_v_b_30')
// (8, 28, 'sp4_v_b_19')
// (8, 29, 'local_g0_6')
// (8, 29, 'ram/RADDR_5')
// (8, 29, 'sp4_h_r_6')
// (8, 29, 'sp4_v_b_6')
// (9, 15, 'sp4_h_r_30')
// (9, 17, 'sp4_h_r_14')
// (9, 21, 'sp12_h_r_4')
// (9, 21, 'sp4_h_r_14')
// (9, 21, 'sp4_h_r_36')
// (9, 29, 'sp4_h_r_19')
// (10, 15, 'sp4_h_r_43')
// (10, 17, 'sp4_h_r_27')
// (10, 21, 'sp12_h_r_7')
// (10, 21, 'sp4_h_l_36')
// (10, 21, 'sp4_h_r_27')
// (10, 29, 'sp4_h_r_30')
// (11, 15, 'sp4_h_l_43')
// (11, 17, 'sp4_h_r_38')
// (11, 21, 'sp12_h_r_8')
// (11, 21, 'sp4_h_r_38')
// (11, 29, 'sp4_h_r_43')
// (12, 17, 'sp4_h_l_38')
// (12, 21, 'sp12_h_r_11')
// (12, 21, 'sp4_h_l_38')
// (12, 29, 'sp4_h_l_43')
// (12, 29, 'sp4_h_r_10')
// (13, 21, 'sp12_h_r_12')
// (13, 29, 'sp4_h_r_23')
// (14, 21, 'sp12_h_r_15')
// (14, 29, 'sp4_h_r_34')
// (15, 21, 'sp12_h_r_16')
// (15, 29, 'sp4_h_r_47')
// (16, 21, 'sp12_h_r_19')
// (16, 29, 'sp4_h_l_47')
// (16, 29, 'sp4_h_r_7')
// (17, 21, 'sp12_h_r_20')
// (17, 29, 'sp4_h_r_18')
// (18, 21, 'sp12_h_r_23')
// (18, 29, 'sp4_h_r_31')
// (19, 18, 'sp4_r_v_b_45')
// (19, 19, 'sp4_r_v_b_32')
// (19, 20, 'sp4_r_v_b_21')
// (19, 21, 'sp12_h_l_23')
// (19, 21, 'sp12_h_r_0')
// (19, 21, 'sp4_r_v_b_8')
// (19, 29, 'sp4_h_r_42')
// (20, 17, 'sp4_v_t_45')
// (20, 18, 'sp4_v_b_45')
// (20, 19, 'local_g2_0')
// (20, 19, 'lutff_7/in_3')
// (20, 19, 'sp4_v_b_32')
// (20, 20, 'sp4_v_b_21')
// (20, 21, 'sp12_h_r_3')
// (20, 21, 'sp4_h_r_3')
// (20, 21, 'sp4_v_b_8')
// (20, 29, 'sp4_h_l_42')
// (20, 29, 'sp4_h_r_4')
// (21, 21, 'sp12_h_r_4')
// (21, 21, 'sp4_h_r_14')
// (21, 29, 'sp4_h_r_17')
// (22, 21, 'sp12_h_r_7')
// (22, 21, 'sp4_h_r_27')
// (22, 29, 'sp4_h_r_28')
// (23, 15, 'sp4_h_r_1')
// (23, 17, 'sp4_h_r_7')
// (23, 19, 'sp4_h_r_4')
// (23, 21, 'local_g1_0')
// (23, 21, 'lutff_0/in_3')
// (23, 21, 'sp12_h_r_8')
// (23, 21, 'sp4_h_r_38')
// (23, 23, 'sp4_h_r_11')
// (23, 29, 'sp4_h_r_41')
// (24, 15, 'sp4_h_r_12')
// (24, 17, 'sp4_h_r_18')
// (24, 19, 'sp4_h_r_17')
// (24, 21, 'sp12_h_r_11')
// (24, 21, 'sp4_h_l_38')
// (24, 23, 'sp4_h_r_22')
// (24, 25, 'sp4_h_r_4')
// (24, 27, 'sp4_h_r_10')
// (24, 29, 'sp4_h_l_41')
// (24, 29, 'sp4_h_r_1')
// (25, 15, 'local_g3_1')
// (25, 15, 'ram/RADDR_5')
// (25, 15, 'sp4_h_r_25')
// (25, 17, 'local_g3_7')
// (25, 17, 'ram/RADDR_5')
// (25, 17, 'sp4_h_r_31')
// (25, 19, 'local_g2_4')
// (25, 19, 'ram/RADDR_5')
// (25, 19, 'sp4_h_r_28')
// (25, 21, 'local_g0_4')
// (25, 21, 'ram/RADDR_5')
// (25, 21, 'sp12_h_r_12')
// (25, 23, 'local_g3_3')
// (25, 23, 'ram/RADDR_5')
// (25, 23, 'sp4_h_r_35')
// (25, 25, 'local_g1_1')
// (25, 25, 'ram/RADDR_5')
// (25, 25, 'sp4_h_r_17')
// (25, 27, 'local_g1_7')
// (25, 27, 'ram/RADDR_5')
// (25, 27, 'sp4_h_r_23')
// (25, 29, 'local_g0_4')
// (25, 29, 'ram/RADDR_5')
// (25, 29, 'sp4_h_r_12')
// (26, 15, 'sp4_h_r_36')
// (26, 17, 'sp4_h_r_42')
// (26, 19, 'sp4_h_r_41')
// (26, 21, 'sp12_h_r_15')
// (26, 23, 'sp4_h_r_46')
// (26, 25, 'sp4_h_r_28')
// (26, 27, 'sp4_h_r_34')
// (26, 29, 'sp4_h_r_25')
// (27, 15, 'sp4_h_l_36')
// (27, 15, 'sp4_h_r_1')
// (27, 17, 'sp4_h_l_42')
// (27, 17, 'sp4_h_r_4')
// (27, 19, 'sp4_h_l_41')
// (27, 19, 'sp4_h_r_4')
// (27, 21, 'sp12_h_r_16')
// (27, 23, 'sp4_h_l_46')
// (27, 23, 'sp4_h_r_3')
// (27, 25, 'sp4_h_r_41')
// (27, 26, 'sp4_r_v_b_41')
// (27, 27, 'sp4_h_r_47')
// (27, 27, 'sp4_r_v_b_28')
// (27, 28, 'sp4_r_v_b_17')
// (27, 28, 'sp4_r_v_b_41')
// (27, 29, 'sp4_h_r_36')
// (27, 29, 'sp4_r_v_b_28')
// (27, 29, 'sp4_r_v_b_4')
// (27, 30, 'sp4_r_v_b_17')
// (27, 30, 'sp4_r_v_b_36')
// (27, 31, 'sp4_r_v_b_25')
// (27, 31, 'sp4_r_v_b_4')
// (27, 32, 'sp4_r_v_b_12')
// (27, 32, 'sp4_r_v_b_36')
// (28, 15, 'sp4_h_r_12')
// (28, 17, 'sp4_h_r_17')
// (28, 19, 'sp4_h_r_17')
// (28, 21, 'sp12_h_r_19')
// (28, 23, 'sp4_h_r_14')
// (28, 25, 'sp4_h_l_41')
// (28, 25, 'sp4_v_t_41')
// (28, 26, 'sp4_v_b_41')
// (28, 27, 'sp4_h_l_47')
// (28, 27, 'sp4_v_b_28')
// (28, 27, 'sp4_v_t_41')
// (28, 28, 'sp4_v_b_17')
// (28, 28, 'sp4_v_b_41')
// (28, 29, 'sp4_h_l_36')
// (28, 29, 'sp4_v_b_28')
// (28, 29, 'sp4_v_b_4')
// (28, 29, 'sp4_v_t_36')
// (28, 30, 'sp4_v_b_17')
// (28, 30, 'sp4_v_b_36')
// (28, 31, 'sp4_v_b_25')
// (28, 31, 'sp4_v_b_4')
// (28, 31, 'sp4_v_t_36')
// (28, 32, 'sp4_v_b_12')
// (28, 32, 'sp4_v_b_36')
// (28, 33, 'span4_horz_r_0')
// (28, 33, 'span4_vert_1')
// (28, 33, 'span4_vert_25')
// (29, 15, 'sp4_h_r_25')
// (29, 17, 'sp4_h_r_28')
// (29, 19, 'sp4_h_r_28')
// (29, 21, 'sp12_h_r_20')
// (29, 23, 'sp4_h_r_27')
// (29, 33, 'span4_horz_r_4')
// (30, 15, 'sp4_h_r_36')
// (30, 16, 'sp4_r_v_b_36')
// (30, 17, 'sp4_h_r_41')
// (30, 17, 'sp4_r_v_b_25')
// (30, 18, 'sp4_r_v_b_12')
// (30, 18, 'sp4_r_v_b_41')
// (30, 19, 'sp4_h_r_41')
// (30, 19, 'sp4_r_v_b_1')
// (30, 19, 'sp4_r_v_b_28')
// (30, 20, 'sp4_r_v_b_17')
// (30, 20, 'sp4_r_v_b_47')
// (30, 21, 'sp12_h_r_23')
// (30, 21, 'sp4_r_v_b_34')
// (30, 21, 'sp4_r_v_b_4')
// (30, 22, 'sp4_r_v_b_23')
// (30, 22, 'sp4_r_v_b_45')
// (30, 23, 'sp4_h_r_38')
// (30, 23, 'sp4_r_v_b_10')
// (30, 23, 'sp4_r_v_b_32')
// (30, 24, 'sp4_r_v_b_21')
// (30, 25, 'sp4_r_v_b_8')
// (30, 32, 'neigh_op_tnr_0')
// (30, 32, 'neigh_op_tnr_4')
// (30, 33, 'span4_horz_r_8')
// (31, 15, 'sp4_h_l_36')
// (31, 15, 'sp4_v_t_36')
// (31, 16, 'sp4_v_b_36')
// (31, 17, 'sp4_h_l_41')
// (31, 17, 'sp4_v_b_25')
// (31, 17, 'sp4_v_t_41')
// (31, 18, 'sp4_v_b_12')
// (31, 18, 'sp4_v_b_41')
// (31, 19, 'sp4_h_l_41')
// (31, 19, 'sp4_v_b_1')
// (31, 19, 'sp4_v_b_28')
// (31, 19, 'sp4_v_t_47')
// (31, 20, 'sp4_v_b_17')
// (31, 20, 'sp4_v_b_47')
// (31, 21, 'sp12_h_l_23')
// (31, 21, 'sp12_v_t_23')
// (31, 21, 'sp4_v_b_34')
// (31, 21, 'sp4_v_b_4')
// (31, 21, 'sp4_v_t_45')
// (31, 22, 'sp12_v_b_23')
// (31, 22, 'sp4_v_b_23')
// (31, 22, 'sp4_v_b_45')
// (31, 23, 'sp12_v_b_20')
// (31, 23, 'sp4_h_l_38')
// (31, 23, 'sp4_v_b_10')
// (31, 23, 'sp4_v_b_32')
// (31, 24, 'sp12_v_b_19')
// (31, 24, 'sp4_v_b_21')
// (31, 25, 'sp12_v_b_16')
// (31, 25, 'sp4_v_b_8')
// (31, 26, 'sp12_v_b_15')
// (31, 27, 'sp12_v_b_12')
// (31, 28, 'sp12_v_b_11')
// (31, 29, 'sp12_v_b_8')
// (31, 30, 'sp12_v_b_7')
// (31, 31, 'sp12_v_b_4')
// (31, 32, 'neigh_op_top_0')
// (31, 32, 'neigh_op_top_4')
// (31, 32, 'sp12_v_b_3')
// (31, 33, 'io_0/D_IN_0')
// (31, 33, 'io_0/PAD')
// (31, 33, 'span12_vert_0')
// (31, 33, 'span4_horz_r_12')
// (32, 32, 'neigh_op_tnl_0')
// (32, 32, 'neigh_op_tnl_4')
// (32, 33, 'span4_horz_l_12')

wire io_31_33_1;
// (6, 12, 'sp4_r_v_b_45')
// (6, 13, 'sp4_r_v_b_32')
// (6, 14, 'sp4_r_v_b_21')
// (6, 14, 'sp4_r_v_b_43')
// (6, 15, 'sp4_r_v_b_30')
// (6, 15, 'sp4_r_v_b_8')
// (6, 16, 'sp4_r_v_b_19')
// (6, 16, 'sp4_r_v_b_41')
// (6, 17, 'sp4_r_v_b_28')
// (6, 17, 'sp4_r_v_b_6')
// (6, 18, 'sp4_r_v_b_17')
// (6, 19, 'sp4_r_v_b_4')
// (7, 11, 'sp12_v_t_23')
// (7, 11, 'sp4_v_t_45')
// (7, 12, 'sp12_v_b_23')
// (7, 12, 'sp4_v_b_45')
// (7, 13, 'sp12_v_b_20')
// (7, 13, 'sp4_v_b_32')
// (7, 13, 'sp4_v_t_43')
// (7, 14, 'sp12_v_b_19')
// (7, 14, 'sp4_v_b_21')
// (7, 14, 'sp4_v_b_43')
// (7, 15, 'sp12_v_b_16')
// (7, 15, 'sp4_h_r_8')
// (7, 15, 'sp4_v_b_30')
// (7, 15, 'sp4_v_b_8')
// (7, 15, 'sp4_v_t_41')
// (7, 16, 'sp12_v_b_15')
// (7, 16, 'sp4_v_b_19')
// (7, 16, 'sp4_v_b_41')
// (7, 17, 'sp12_v_b_12')
// (7, 17, 'sp4_h_r_0')
// (7, 17, 'sp4_v_b_28')
// (7, 17, 'sp4_v_b_6')
// (7, 18, 'sp12_v_b_11')
// (7, 18, 'sp4_v_b_17')
// (7, 19, 'sp12_v_b_8')
// (7, 19, 'sp4_h_r_4')
// (7, 19, 'sp4_v_b_4')
// (7, 20, 'sp12_v_b_7')
// (7, 20, 'sp4_r_v_b_38')
// (7, 21, 'sp12_v_b_4')
// (7, 21, 'sp4_r_v_b_27')
// (7, 22, 'sp12_v_b_3')
// (7, 22, 'sp4_r_v_b_14')
// (7, 23, 'sp12_h_r_0')
// (7, 23, 'sp12_v_b_0')
// (7, 23, 'sp4_r_v_b_3')
// (7, 24, 'sp4_r_v_b_44')
// (7, 25, 'sp4_r_v_b_33')
// (7, 26, 'sp4_r_v_b_20')
// (7, 27, 'sp12_h_r_0')
// (7, 27, 'sp4_r_v_b_9')
// (7, 29, 'sp4_h_r_3')
// (8, 15, 'local_g0_5')
// (8, 15, 'ram/RADDR_4')
// (8, 15, 'sp4_h_r_21')
// (8, 17, 'local_g0_5')
// (8, 17, 'ram/RADDR_4')
// (8, 17, 'sp4_h_r_13')
// (8, 19, 'local_g0_1')
// (8, 19, 'ram/RADDR_4')
// (8, 19, 'sp4_h_r_17')
// (8, 19, 'sp4_v_t_38')
// (8, 20, 'sp4_v_b_38')
// (8, 21, 'local_g2_3')
// (8, 21, 'ram/RADDR_4')
// (8, 21, 'sp4_v_b_27')
// (8, 22, 'sp4_v_b_14')
// (8, 23, 'local_g0_3')
// (8, 23, 'ram/RADDR_4')
// (8, 23, 'sp12_h_r_3')
// (8, 23, 'sp4_h_r_3')
// (8, 23, 'sp4_v_b_3')
// (8, 23, 'sp4_v_t_44')
// (8, 24, 'sp4_v_b_44')
// (8, 25, 'local_g2_1')
// (8, 25, 'ram/RADDR_4')
// (8, 25, 'sp4_v_b_33')
// (8, 26, 'sp4_v_b_20')
// (8, 27, 'local_g0_3')
// (8, 27, 'ram/RADDR_4')
// (8, 27, 'sp12_h_r_3')
// (8, 27, 'sp4_v_b_9')
// (8, 29, 'local_g1_6')
// (8, 29, 'ram/RADDR_4')
// (8, 29, 'sp4_h_r_14')
// (9, 15, 'sp4_h_r_32')
// (9, 17, 'sp4_h_r_24')
// (9, 19, 'sp4_h_r_28')
// (9, 23, 'sp12_h_r_4')
// (9, 23, 'sp4_h_r_14')
// (9, 27, 'sp12_h_r_4')
// (9, 29, 'sp4_h_r_27')
// (10, 15, 'sp4_h_r_45')
// (10, 17, 'sp4_h_r_37')
// (10, 19, 'sp4_h_r_41')
// (10, 23, 'sp12_h_r_7')
// (10, 23, 'sp4_h_r_27')
// (10, 27, 'sp12_h_r_7')
// (10, 29, 'sp4_h_r_38')
// (11, 15, 'sp4_h_l_45')
// (11, 17, 'sp4_h_l_37')
// (11, 19, 'sp4_h_l_41')
// (11, 23, 'sp12_h_r_8')
// (11, 23, 'sp4_h_r_38')
// (11, 27, 'sp12_h_r_8')
// (11, 29, 'sp4_h_l_38')
// (11, 29, 'sp4_h_r_0')
// (12, 23, 'sp12_h_r_11')
// (12, 23, 'sp4_h_l_38')
// (12, 27, 'sp12_h_r_11')
// (12, 29, 'sp4_h_r_13')
// (13, 23, 'sp12_h_r_12')
// (13, 27, 'sp12_h_r_12')
// (13, 29, 'sp4_h_r_24')
// (14, 23, 'sp12_h_r_15')
// (14, 27, 'sp12_h_r_15')
// (14, 29, 'sp4_h_r_37')
// (15, 23, 'sp12_h_r_16')
// (15, 27, 'sp12_h_r_16')
// (15, 29, 'sp4_h_l_37')
// (15, 29, 'sp4_h_r_4')
// (16, 23, 'sp12_h_r_19')
// (16, 27, 'sp12_h_r_19')
// (16, 29, 'sp4_h_r_17')
// (17, 23, 'sp12_h_r_20')
// (17, 27, 'sp12_h_r_20')
// (17, 29, 'sp4_h_r_28')
// (18, 23, 'sp12_h_r_23')
// (18, 27, 'sp12_h_r_23')
// (18, 29, 'sp4_h_r_41')
// (19, 15, 'sp12_h_r_0')
// (19, 20, 'sp4_r_v_b_38')
// (19, 21, 'sp4_r_v_b_27')
// (19, 22, 'sp4_r_v_b_14')
// (19, 23, 'sp12_h_l_23')
// (19, 23, 'sp12_h_r_0')
// (19, 23, 'sp4_r_v_b_3')
// (19, 27, 'sp12_h_l_23')
// (19, 27, 'sp12_h_r_0')
// (19, 29, 'sp4_h_l_41')
// (19, 29, 'sp4_h_r_8')
// (20, 15, 'sp12_h_r_3')
// (20, 19, 'local_g0_0')
// (20, 19, 'lutff_6/in_2')
// (20, 19, 'sp4_h_r_8')
// (20, 19, 'sp4_v_t_38')
// (20, 20, 'sp4_v_b_38')
// (20, 21, 'sp4_v_b_27')
// (20, 22, 'sp4_v_b_14')
// (20, 23, 'sp12_h_r_3')
// (20, 23, 'sp4_h_r_3')
// (20, 23, 'sp4_v_b_3')
// (20, 27, 'sp12_h_r_3')
// (20, 29, 'sp4_h_r_21')
// (21, 15, 'sp12_h_r_4')
// (21, 19, 'sp4_h_r_21')
// (21, 23, 'sp12_h_r_4')
// (21, 23, 'sp4_h_r_14')
// (21, 27, 'sp12_h_r_4')
// (21, 29, 'sp4_h_r_32')
// (22, 15, 'sp12_h_r_7')
// (22, 19, 'sp4_h_r_32')
// (22, 23, 'sp12_h_r_7')
// (22, 23, 'sp4_h_r_27')
// (22, 23, 'sp4_h_r_5')
// (22, 27, 'sp12_h_r_7')
// (22, 29, 'sp4_h_r_45')
// (23, 15, 'sp12_h_r_8')
// (23, 17, 'sp4_h_r_3')
// (23, 19, 'sp4_h_r_45')
// (23, 20, 'sp4_r_v_b_38')
// (23, 21, 'local_g1_6')
// (23, 21, 'lutff_0/in_1')
// (23, 21, 'sp4_h_r_6')
// (23, 21, 'sp4_r_v_b_27')
// (23, 22, 'sp4_r_v_b_14')
// (23, 23, 'sp12_h_r_8')
// (23, 23, 'sp4_h_r_16')
// (23, 23, 'sp4_h_r_38')
// (23, 23, 'sp4_r_v_b_3')
// (23, 25, 'sp4_h_r_0')
// (23, 27, 'sp12_h_r_8')
// (23, 29, 'sp4_h_l_45')
// (23, 29, 'sp4_h_r_0')
// (24, 15, 'sp12_h_r_11')
// (24, 17, 'sp4_h_r_14')
// (24, 19, 'sp4_h_l_45')
// (24, 19, 'sp4_h_r_8')
// (24, 19, 'sp4_v_t_38')
// (24, 20, 'sp4_v_b_38')
// (24, 21, 'sp4_h_r_19')
// (24, 21, 'sp4_v_b_27')
// (24, 22, 'sp4_v_b_14')
// (24, 23, 'sp12_h_r_11')
// (24, 23, 'sp4_h_l_38')
// (24, 23, 'sp4_h_r_29')
// (24, 23, 'sp4_v_b_3')
// (24, 25, 'sp4_h_r_13')
// (24, 27, 'sp12_h_r_11')
// (24, 27, 'sp4_h_r_7')
// (24, 29, 'sp4_h_r_13')
// (25, 15, 'local_g1_4')
// (25, 15, 'ram/RADDR_4')
// (25, 15, 'sp12_h_r_12')
// (25, 17, 'local_g2_3')
// (25, 17, 'ram/RADDR_4')
// (25, 17, 'sp4_h_r_27')
// (25, 19, 'local_g0_5')
// (25, 19, 'ram/RADDR_4')
// (25, 19, 'sp4_h_r_21')
// (25, 21, 'local_g3_6')
// (25, 21, 'ram/RADDR_4')
// (25, 21, 'sp4_h_r_30')
// (25, 23, 'local_g3_0')
// (25, 23, 'ram/RADDR_4')
// (25, 23, 'sp12_h_r_12')
// (25, 23, 'sp4_h_r_40')
// (25, 25, 'local_g3_0')
// (25, 25, 'ram/RADDR_4')
// (25, 25, 'sp4_h_r_24')
// (25, 27, 'local_g1_2')
// (25, 27, 'ram/RADDR_4')
// (25, 27, 'sp12_h_r_12')
// (25, 27, 'sp4_h_r_18')
// (25, 29, 'local_g3_0')
// (25, 29, 'ram/RADDR_4')
// (25, 29, 'sp4_h_r_24')
// (26, 15, 'sp12_h_r_15')
// (26, 17, 'sp4_h_r_38')
// (26, 18, 'sp4_r_v_b_38')
// (26, 19, 'sp4_h_r_32')
// (26, 19, 'sp4_r_v_b_27')
// (26, 20, 'sp4_r_v_b_14')
// (26, 21, 'sp4_h_r_43')
// (26, 21, 'sp4_r_v_b_3')
// (26, 23, 'sp12_h_r_15')
// (26, 23, 'sp4_h_l_40')
// (26, 25, 'sp4_h_r_37')
// (26, 27, 'sp12_h_r_15')
// (26, 27, 'sp4_h_r_31')
// (26, 29, 'sp4_h_r_37')
// (27, 15, 'sp12_h_r_16')
// (27, 17, 'sp4_h_l_38')
// (27, 17, 'sp4_v_t_38')
// (27, 18, 'sp4_v_b_38')
// (27, 19, 'sp4_h_r_45')
// (27, 19, 'sp4_v_b_27')
// (27, 20, 'sp4_v_b_14')
// (27, 21, 'sp4_h_l_43')
// (27, 21, 'sp4_h_r_10')
// (27, 21, 'sp4_v_b_3')
// (27, 23, 'sp12_h_r_16')
// (27, 25, 'sp4_h_l_37')
// (27, 25, 'sp4_h_r_0')
// (27, 27, 'sp12_h_r_16')
// (27, 27, 'sp4_h_r_42')
// (27, 29, 'sp4_h_l_37')
// (27, 29, 'sp4_h_r_4')
// (28, 15, 'sp12_h_r_19')
// (28, 19, 'sp4_h_l_45')
// (28, 21, 'sp4_h_r_23')
// (28, 23, 'sp12_h_r_19')
// (28, 25, 'sp4_h_r_13')
// (28, 27, 'sp12_h_r_19')
// (28, 27, 'sp4_h_l_42')
// (28, 29, 'sp4_h_r_17')
// (29, 15, 'sp12_h_r_20')
// (29, 21, 'sp4_h_r_34')
// (29, 23, 'sp12_h_r_20')
// (29, 25, 'sp4_h_r_24')
// (29, 27, 'sp12_h_r_20')
// (29, 29, 'sp4_h_r_28')
// (30, 15, 'sp12_h_r_23')
// (30, 21, 'sp4_h_r_47')
// (30, 22, 'sp4_r_v_b_47')
// (30, 23, 'sp12_h_r_23')
// (30, 23, 'sp4_r_v_b_34')
// (30, 24, 'sp4_r_v_b_23')
// (30, 25, 'sp4_h_r_37')
// (30, 25, 'sp4_r_v_b_10')
// (30, 26, 'sp4_r_v_b_37')
// (30, 27, 'sp12_h_r_23')
// (30, 27, 'sp4_r_v_b_24')
// (30, 28, 'sp4_r_v_b_13')
// (30, 29, 'sp4_h_r_41')
// (30, 29, 'sp4_r_v_b_0')
// (30, 30, 'sp4_r_v_b_41')
// (30, 31, 'sp4_r_v_b_28')
// (30, 32, 'neigh_op_tnr_2')
// (30, 32, 'neigh_op_tnr_6')
// (30, 32, 'sp4_r_v_b_17')
// (31, 15, 'sp12_h_l_23')
// (31, 15, 'sp12_v_t_23')
// (31, 16, 'sp12_v_b_23')
// (31, 17, 'sp12_v_b_20')
// (31, 18, 'sp12_v_b_19')
// (31, 19, 'sp12_v_b_16')
// (31, 20, 'sp12_v_b_15')
// (31, 21, 'sp12_v_b_12')
// (31, 21, 'sp4_h_l_47')
// (31, 21, 'sp4_v_t_47')
// (31, 22, 'sp12_v_b_11')
// (31, 22, 'sp4_v_b_47')
// (31, 23, 'sp12_h_l_23')
// (31, 23, 'sp12_v_b_8')
// (31, 23, 'sp12_v_t_23')
// (31, 23, 'sp4_v_b_34')
// (31, 24, 'sp12_v_b_23')
// (31, 24, 'sp12_v_b_7')
// (31, 24, 'sp4_v_b_23')
// (31, 25, 'sp12_v_b_20')
// (31, 25, 'sp12_v_b_4')
// (31, 25, 'sp4_h_l_37')
// (31, 25, 'sp4_v_b_10')
// (31, 25, 'sp4_v_t_37')
// (31, 26, 'sp12_v_b_19')
// (31, 26, 'sp12_v_b_3')
// (31, 26, 'sp4_v_b_37')
// (31, 27, 'sp12_h_l_23')
// (31, 27, 'sp12_v_b_0')
// (31, 27, 'sp12_v_b_16')
// (31, 27, 'sp12_v_t_23')
// (31, 27, 'sp4_v_b_24')
// (31, 28, 'sp12_v_b_15')
// (31, 28, 'sp12_v_b_23')
// (31, 28, 'sp4_v_b_13')
// (31, 29, 'sp12_v_b_12')
// (31, 29, 'sp12_v_b_20')
// (31, 29, 'sp4_h_l_41')
// (31, 29, 'sp4_v_b_0')
// (31, 29, 'sp4_v_t_41')
// (31, 30, 'sp12_v_b_11')
// (31, 30, 'sp12_v_b_19')
// (31, 30, 'sp4_v_b_41')
// (31, 31, 'sp12_v_b_16')
// (31, 31, 'sp12_v_b_8')
// (31, 31, 'sp4_v_b_28')
// (31, 32, 'neigh_op_top_2')
// (31, 32, 'neigh_op_top_6')
// (31, 32, 'sp12_v_b_15')
// (31, 32, 'sp12_v_b_7')
// (31, 32, 'sp4_v_b_17')
// (31, 33, 'io_1/D_IN_0')
// (31, 33, 'io_1/PAD')
// (31, 33, 'span12_vert_12')
// (31, 33, 'span12_vert_4')
// (31, 33, 'span4_vert_4')
// (32, 32, 'neigh_op_tnl_2')
// (32, 32, 'neigh_op_tnl_6')

wire n36;
// (6, 16, 'sp4_r_v_b_45')
// (6, 17, 'sp4_r_v_b_32')
// (6, 18, 'neigh_op_tnr_4')
// (6, 18, 'sp4_r_v_b_21')
// (6, 19, 'neigh_op_rgt_4')
// (6, 19, 'sp4_r_v_b_8')
// (6, 20, 'neigh_op_bnr_4')
// (7, 15, 'sp4_v_t_45')
// (7, 16, 'sp4_v_b_45')
// (7, 17, 'sp4_v_b_32')
// (7, 18, 'neigh_op_top_4')
// (7, 18, 'sp4_v_b_21')
// (7, 19, 'local_g0_0')
// (7, 19, 'lutff_0/in_0')
// (7, 19, 'lutff_4/out')
// (7, 19, 'sp4_v_b_8')
// (7, 20, 'neigh_op_bot_4')
// (8, 18, 'neigh_op_tnl_4')
// (8, 19, 'neigh_op_lft_4')
// (8, 20, 'neigh_op_bnl_4')

wire n37;
// (6, 18, 'neigh_op_tnr_2')
// (6, 19, 'neigh_op_rgt_2')
// (6, 20, 'neigh_op_bnr_2')
// (7, 18, 'neigh_op_top_2')
// (7, 19, 'local_g3_2')
// (7, 19, 'lutff_2/out')
// (7, 19, 'lutff_3/in_2')
// (7, 20, 'neigh_op_bot_2')
// (8, 18, 'neigh_op_tnl_2')
// (8, 19, 'neigh_op_lft_2')
// (8, 20, 'neigh_op_bnl_2')

reg n38 = 0;
// (6, 19, 'neigh_op_tnr_2')
// (6, 20, 'neigh_op_rgt_2')
// (6, 21, 'neigh_op_bnr_2')
// (7, 19, 'neigh_op_top_2')
// (7, 20, 'local_g2_2')
// (7, 20, 'lutff_2/in_2')
// (7, 20, 'lutff_2/out')
// (7, 20, 'sp4_r_v_b_37')
// (7, 21, 'neigh_op_bot_2')
// (7, 21, 'sp4_r_v_b_24')
// (7, 22, 'local_g2_5')
// (7, 22, 'lutff_5/in_2')
// (7, 22, 'sp4_r_v_b_13')
// (7, 23, 'sp4_r_v_b_0')
// (8, 19, 'neigh_op_tnl_2')
// (8, 19, 'sp4_v_t_37')
// (8, 20, 'neigh_op_lft_2')
// (8, 20, 'sp4_v_b_37')
// (8, 21, 'neigh_op_bnl_2')
// (8, 21, 'sp4_v_b_24')
// (8, 22, 'sp4_v_b_13')
// (8, 23, 'sp4_v_b_0')

reg n39 = 0;
// (6, 19, 'neigh_op_tnr_3')
// (6, 20, 'neigh_op_rgt_3')
// (6, 21, 'neigh_op_bnr_3')
// (7, 19, 'neigh_op_top_3')
// (7, 20, 'local_g2_3')
// (7, 20, 'lutff_3/in_2')
// (7, 20, 'lutff_3/out')
// (7, 21, 'local_g0_3')
// (7, 21, 'lutff_4/in_3')
// (7, 21, 'neigh_op_bot_3')
// (8, 19, 'neigh_op_tnl_3')
// (8, 20, 'neigh_op_lft_3')
// (8, 21, 'neigh_op_bnl_3')

reg n40 = 0;
// (6, 19, 'neigh_op_tnr_4')
// (6, 20, 'neigh_op_rgt_4')
// (6, 21, 'neigh_op_bnr_4')
// (7, 19, 'local_g1_4')
// (7, 19, 'lutff_0/in_1')
// (7, 19, 'neigh_op_top_4')
// (7, 20, 'local_g0_4')
// (7, 20, 'lutff_4/in_2')
// (7, 20, 'lutff_4/out')
// (7, 21, 'neigh_op_bot_4')
// (8, 19, 'neigh_op_tnl_4')
// (8, 20, 'neigh_op_lft_4')
// (8, 21, 'neigh_op_bnl_4')

reg n41 = 0;
// (6, 19, 'neigh_op_tnr_5')
// (6, 20, 'neigh_op_rgt_5')
// (6, 21, 'neigh_op_bnr_5')
// (7, 19, 'local_g1_5')
// (7, 19, 'lutff_3/in_3')
// (7, 19, 'neigh_op_top_5')
// (7, 20, 'local_g1_5')
// (7, 20, 'lutff_5/in_1')
// (7, 20, 'lutff_5/out')
// (7, 21, 'neigh_op_bot_5')
// (8, 19, 'neigh_op_tnl_5')
// (8, 20, 'neigh_op_lft_5')
// (8, 21, 'neigh_op_bnl_5')

reg n42 = 0;
// (6, 19, 'neigh_op_tnr_6')
// (6, 20, 'neigh_op_rgt_6')
// (6, 21, 'neigh_op_bnr_6')
// (7, 19, 'neigh_op_top_6')
// (7, 20, 'local_g1_6')
// (7, 20, 'lutff_6/in_1')
// (7, 20, 'lutff_6/out')
// (7, 21, 'local_g0_6')
// (7, 21, 'lutff_7/in_3')
// (7, 21, 'neigh_op_bot_6')
// (8, 19, 'neigh_op_tnl_6')
// (8, 20, 'neigh_op_lft_6')
// (8, 21, 'neigh_op_bnl_6')

reg n43 = 0;
// (6, 19, 'neigh_op_tnr_7')
// (6, 20, 'neigh_op_rgt_7')
// (6, 21, 'neigh_op_bnr_7')
// (7, 19, 'neigh_op_top_7')
// (7, 20, 'local_g2_7')
// (7, 20, 'lutff_7/in_2')
// (7, 20, 'lutff_7/out')
// (7, 21, 'local_g1_7')
// (7, 21, 'lutff_5/in_3')
// (7, 21, 'neigh_op_bot_7')
// (8, 19, 'neigh_op_tnl_7')
// (8, 20, 'neigh_op_lft_7')
// (8, 21, 'neigh_op_bnl_7')

wire n44;
// (6, 20, 'neigh_op_tnr_2')
// (6, 21, 'neigh_op_rgt_2')
// (6, 22, 'neigh_op_bnr_2')
// (7, 20, 'neigh_op_top_2')
// (7, 21, 'local_g0_2')
// (7, 21, 'lutff_2/out')
// (7, 21, 'lutff_7/in_1')
// (7, 22, 'neigh_op_bot_2')
// (8, 20, 'neigh_op_tnl_2')
// (8, 21, 'neigh_op_lft_2')
// (8, 22, 'neigh_op_bnl_2')

wire n45;
// (6, 20, 'neigh_op_tnr_6')
// (6, 21, 'neigh_op_rgt_6')
// (6, 22, 'neigh_op_bnr_6')
// (7, 20, 'neigh_op_top_6')
// (7, 21, 'local_g2_6')
// (7, 21, 'lutff_5/in_1')
// (7, 21, 'lutff_6/out')
// (7, 22, 'neigh_op_bot_6')
// (8, 20, 'neigh_op_tnl_6')
// (8, 21, 'neigh_op_lft_6')
// (8, 22, 'neigh_op_bnl_6')

wire n46;
// (6, 20, 'sp4_r_v_b_37')
// (6, 21, 'sp4_r_v_b_24')
// (6, 22, 'neigh_op_tnr_0')
// (6, 22, 'sp4_r_v_b_13')
// (6, 23, 'neigh_op_rgt_0')
// (6, 23, 'sp4_r_v_b_0')
// (6, 24, 'neigh_op_bnr_0')
// (7, 19, 'sp4_v_t_37')
// (7, 20, 'sp4_v_b_37')
// (7, 21, 'local_g2_0')
// (7, 21, 'lutff_1/in_1')
// (7, 21, 'sp4_v_b_24')
// (7, 22, 'neigh_op_top_0')
// (7, 22, 'sp4_v_b_13')
// (7, 23, 'lutff_0/out')
// (7, 23, 'sp4_v_b_0')
// (7, 24, 'neigh_op_bot_0')
// (8, 22, 'neigh_op_tnl_0')
// (8, 23, 'neigh_op_lft_0')
// (8, 24, 'neigh_op_bnl_0')

wire io_30_33_0;
// (6, 21, 'sp12_h_r_0')
// (6, 29, 'sp12_h_r_0')
// (7, 21, 'sp12_h_r_3')
// (7, 29, 'sp12_h_r_3')
// (8, 14, 'sp4_r_v_b_40')
// (8, 14, 'sp4_r_v_b_45')
// (8, 15, 'local_g1_5')
// (8, 15, 'ram/RADDR_3')
// (8, 15, 'sp4_r_v_b_29')
// (8, 15, 'sp4_r_v_b_32')
// (8, 16, 'sp4_r_v_b_16')
// (8, 16, 'sp4_r_v_b_21')
// (8, 17, 'local_g2_0')
// (8, 17, 'ram/RADDR_3')
// (8, 17, 'sp4_r_v_b_5')
// (8, 17, 'sp4_r_v_b_8')
// (8, 18, 'sp4_r_v_b_40')
// (8, 19, 'local_g1_5')
// (8, 19, 'ram/RADDR_3')
// (8, 19, 'sp4_r_v_b_29')
// (8, 20, 'sp4_r_v_b_16')
// (8, 21, 'local_g0_4')
// (8, 21, 'ram/RADDR_3')
// (8, 21, 'sp12_h_r_4')
// (8, 21, 'sp4_r_v_b_5')
// (8, 22, 'sp4_r_v_b_40')
// (8, 22, 'sp4_r_v_b_47')
// (8, 23, 'local_g1_5')
// (8, 23, 'ram/RADDR_3')
// (8, 23, 'sp4_r_v_b_29')
// (8, 23, 'sp4_r_v_b_34')
// (8, 24, 'sp4_r_v_b_16')
// (8, 24, 'sp4_r_v_b_23')
// (8, 25, 'local_g2_2')
// (8, 25, 'ram/RADDR_3')
// (8, 25, 'sp4_r_v_b_10')
// (8, 25, 'sp4_r_v_b_5')
// (8, 26, 'sp4_r_v_b_47')
// (8, 27, 'local_g2_2')
// (8, 27, 'ram/RADDR_3')
// (8, 27, 'sp4_r_v_b_34')
// (8, 28, 'sp4_r_v_b_23')
// (8, 29, 'local_g0_4')
// (8, 29, 'ram/RADDR_3')
// (8, 29, 'sp12_h_r_4')
// (8, 29, 'sp4_r_v_b_10')
// (9, 13, 'sp4_v_t_40')
// (9, 13, 'sp4_v_t_45')
// (9, 14, 'sp4_v_b_40')
// (9, 14, 'sp4_v_b_45')
// (9, 15, 'sp4_v_b_29')
// (9, 15, 'sp4_v_b_32')
// (9, 16, 'sp4_v_b_16')
// (9, 16, 'sp4_v_b_21')
// (9, 17, 'sp4_v_b_5')
// (9, 17, 'sp4_v_b_8')
// (9, 17, 'sp4_v_t_40')
// (9, 18, 'sp4_v_b_40')
// (9, 19, 'sp4_v_b_29')
// (9, 20, 'sp4_v_b_16')
// (9, 21, 'sp12_h_r_7')
// (9, 21, 'sp4_h_r_5')
// (9, 21, 'sp4_v_b_5')
// (9, 21, 'sp4_v_t_40')
// (9, 21, 'sp4_v_t_47')
// (9, 22, 'sp4_v_b_40')
// (9, 22, 'sp4_v_b_47')
// (9, 23, 'sp4_v_b_29')
// (9, 23, 'sp4_v_b_34')
// (9, 24, 'sp4_v_b_16')
// (9, 24, 'sp4_v_b_23')
// (9, 25, 'sp4_v_b_10')
// (9, 25, 'sp4_v_b_5')
// (9, 25, 'sp4_v_t_47')
// (9, 26, 'sp4_v_b_47')
// (9, 27, 'sp4_v_b_34')
// (9, 28, 'sp4_v_b_23')
// (9, 29, 'sp12_h_r_7')
// (9, 29, 'sp4_h_r_5')
// (9, 29, 'sp4_v_b_10')
// (10, 21, 'sp12_h_r_8')
// (10, 21, 'sp4_h_r_16')
// (10, 29, 'sp12_h_r_8')
// (10, 29, 'sp4_h_r_16')
// (11, 21, 'sp12_h_r_11')
// (11, 21, 'sp4_h_r_29')
// (11, 29, 'sp12_h_r_11')
// (11, 29, 'sp4_h_r_29')
// (12, 21, 'sp12_h_r_12')
// (12, 21, 'sp4_h_r_40')
// (12, 29, 'sp12_h_r_12')
// (12, 29, 'sp4_h_r_40')
// (13, 21, 'sp12_h_r_15')
// (13, 21, 'sp4_h_l_40')
// (13, 29, 'sp12_h_r_15')
// (13, 29, 'sp4_h_l_40')
// (14, 21, 'sp12_h_r_16')
// (14, 29, 'sp12_h_r_16')
// (15, 21, 'sp12_h_r_19')
// (15, 29, 'sp12_h_r_19')
// (16, 21, 'sp12_h_r_20')
// (16, 29, 'sp12_h_r_20')
// (17, 21, 'sp12_h_r_23')
// (17, 29, 'sp12_h_r_23')
// (18, 21, 'sp12_h_l_23')
// (18, 21, 'sp12_h_r_0')
// (18, 29, 'sp12_h_l_23')
// (18, 29, 'sp12_h_r_0')
// (19, 21, 'sp12_h_r_3')
// (19, 29, 'sp12_h_r_3')
// (20, 21, 'sp12_h_r_4')
// (20, 29, 'sp12_h_r_4')
// (21, 16, 'sp4_r_v_b_40')
// (21, 17, 'sp4_r_v_b_29')
// (21, 18, 'sp4_r_v_b_16')
// (21, 19, 'sp4_r_v_b_5')
// (21, 21, 'sp12_h_r_7')
// (21, 29, 'sp12_h_r_7')
// (22, 15, 'sp4_v_t_40')
// (22, 16, 'sp4_v_b_40')
// (22, 17, 'sp4_v_b_29')
// (22, 18, 'local_g0_0')
// (22, 18, 'lutff_2/in_2')
// (22, 18, 'sp4_v_b_16')
// (22, 19, 'sp4_h_r_0')
// (22, 19, 'sp4_v_b_5')
// (22, 21, 'sp12_h_r_8')
// (22, 29, 'sp12_h_r_8')
// (23, 19, 'sp4_h_r_13')
// (23, 21, 'local_g0_3')
// (23, 21, 'lutff_6/in_3')
// (23, 21, 'sp12_h_r_11')
// (23, 29, 'sp12_h_r_11')
// (24, 19, 'sp4_h_r_24')
// (24, 21, 'sp12_h_r_12')
// (24, 29, 'sp12_h_r_12')
// (25, 12, 'sp4_r_v_b_40')
// (25, 13, 'sp4_r_v_b_29')
// (25, 14, 'sp4_r_v_b_16')
// (25, 15, 'local_g1_5')
// (25, 15, 'ram/RADDR_3')
// (25, 15, 'sp4_r_v_b_5')
// (25, 16, 'sp4_r_v_b_41')
// (25, 16, 'sp4_r_v_b_44')
// (25, 16, 'sp4_r_v_b_47')
// (25, 17, 'local_g0_4')
// (25, 17, 'ram/RADDR_3')
// (25, 17, 'sp4_r_v_b_28')
// (25, 17, 'sp4_r_v_b_33')
// (25, 17, 'sp4_r_v_b_34')
// (25, 18, 'sp4_r_v_b_17')
// (25, 18, 'sp4_r_v_b_20')
// (25, 18, 'sp4_r_v_b_23')
// (25, 19, 'local_g2_2')
// (25, 19, 'ram/RADDR_3')
// (25, 19, 'sp4_h_r_37')
// (25, 19, 'sp4_r_v_b_10')
// (25, 19, 'sp4_r_v_b_4')
// (25, 19, 'sp4_r_v_b_9')
// (25, 20, 'sp4_r_v_b_45')
// (25, 21, 'local_g1_7')
// (25, 21, 'ram/RADDR_3')
// (25, 21, 'sp12_h_r_15')
// (25, 21, 'sp4_r_v_b_32')
// (25, 22, 'sp4_r_v_b_21')
// (25, 22, 'sp4_r_v_b_45')
// (25, 23, 'local_g2_0')
// (25, 23, 'ram/RADDR_3')
// (25, 23, 'sp4_r_v_b_32')
// (25, 23, 'sp4_r_v_b_8')
// (25, 24, 'sp4_r_v_b_21')
// (25, 25, 'local_g2_0')
// (25, 25, 'ram/RADDR_3')
// (25, 25, 'sp4_r_v_b_8')
// (25, 26, 'sp4_r_v_b_36')
// (25, 26, 'sp4_r_v_b_45')
// (25, 27, 'local_g2_0')
// (25, 27, 'ram/RADDR_3')
// (25, 27, 'sp4_r_v_b_25')
// (25, 27, 'sp4_r_v_b_32')
// (25, 28, 'sp4_r_v_b_12')
// (25, 28, 'sp4_r_v_b_21')
// (25, 29, 'local_g1_1')
// (25, 29, 'ram/RADDR_3')
// (25, 29, 'sp12_h_r_15')
// (25, 29, 'sp4_r_v_b_1')
// (25, 29, 'sp4_r_v_b_8')
// (26, 11, 'sp4_v_t_40')
// (26, 12, 'sp4_v_b_40')
// (26, 13, 'sp4_v_b_29')
// (26, 14, 'sp4_v_b_16')
// (26, 15, 'sp4_v_b_5')
// (26, 15, 'sp4_v_t_41')
// (26, 15, 'sp4_v_t_44')
// (26, 15, 'sp4_v_t_47')
// (26, 16, 'sp4_v_b_41')
// (26, 16, 'sp4_v_b_44')
// (26, 16, 'sp4_v_b_47')
// (26, 17, 'sp4_v_b_28')
// (26, 17, 'sp4_v_b_33')
// (26, 17, 'sp4_v_b_34')
// (26, 18, 'sp4_v_b_17')
// (26, 18, 'sp4_v_b_20')
// (26, 18, 'sp4_v_b_23')
// (26, 19, 'sp4_h_l_37')
// (26, 19, 'sp4_h_r_10')
// (26, 19, 'sp4_h_r_4')
// (26, 19, 'sp4_v_b_10')
// (26, 19, 'sp4_v_b_4')
// (26, 19, 'sp4_v_b_9')
// (26, 19, 'sp4_v_t_45')
// (26, 20, 'sp4_v_b_45')
// (26, 21, 'sp12_h_r_16')
// (26, 21, 'sp4_v_b_32')
// (26, 21, 'sp4_v_t_45')
// (26, 22, 'sp4_v_b_21')
// (26, 22, 'sp4_v_b_45')
// (26, 23, 'sp4_h_r_3')
// (26, 23, 'sp4_v_b_32')
// (26, 23, 'sp4_v_b_8')
// (26, 24, 'sp4_v_b_21')
// (26, 25, 'sp4_h_r_8')
// (26, 25, 'sp4_v_b_8')
// (26, 25, 'sp4_v_t_36')
// (26, 25, 'sp4_v_t_45')
// (26, 26, 'sp4_v_b_36')
// (26, 26, 'sp4_v_b_45')
// (26, 27, 'sp4_v_b_25')
// (26, 27, 'sp4_v_b_32')
// (26, 28, 'sp4_v_b_12')
// (26, 28, 'sp4_v_b_21')
// (26, 29, 'sp12_h_r_16')
// (26, 29, 'sp4_h_r_8')
// (26, 29, 'sp4_v_b_1')
// (26, 29, 'sp4_v_b_8')
// (27, 19, 'sp4_h_r_17')
// (27, 19, 'sp4_h_r_23')
// (27, 21, 'sp12_h_r_19')
// (27, 23, 'sp4_h_r_14')
// (27, 25, 'sp4_h_r_21')
// (27, 29, 'sp12_h_r_19')
// (27, 29, 'sp4_h_r_21')
// (28, 19, 'sp4_h_r_28')
// (28, 19, 'sp4_h_r_34')
// (28, 21, 'sp12_h_r_20')
// (28, 23, 'sp4_h_r_27')
// (28, 25, 'sp4_h_r_32')
// (28, 29, 'sp12_h_r_20')
// (28, 29, 'sp4_h_r_32')
// (29, 19, 'sp4_h_r_41')
// (29, 19, 'sp4_h_r_47')
// (29, 20, 'sp4_r_v_b_47')
// (29, 21, 'sp12_h_r_23')
// (29, 21, 'sp4_r_v_b_34')
// (29, 22, 'sp4_r_v_b_23')
// (29, 23, 'sp4_h_r_38')
// (29, 23, 'sp4_r_v_b_10')
// (29, 25, 'sp4_h_r_45')
// (29, 26, 'sp4_r_v_b_45')
// (29, 27, 'sp4_r_v_b_32')
// (29, 28, 'sp4_r_v_b_21')
// (29, 29, 'sp12_h_r_23')
// (29, 29, 'sp4_h_r_45')
// (29, 29, 'sp4_r_v_b_8')
// (29, 30, 'sp4_r_v_b_45')
// (29, 31, 'sp4_r_v_b_32')
// (29, 32, 'neigh_op_tnr_0')
// (29, 32, 'neigh_op_tnr_4')
// (29, 32, 'sp4_r_v_b_21')
// (30, 19, 'sp4_h_l_41')
// (30, 19, 'sp4_h_l_47')
// (30, 19, 'sp4_v_t_47')
// (30, 20, 'sp4_v_b_47')
// (30, 21, 'sp12_h_l_23')
// (30, 21, 'sp12_v_t_23')
// (30, 21, 'sp4_v_b_34')
// (30, 22, 'sp12_v_b_23')
// (30, 22, 'sp4_v_b_23')
// (30, 23, 'sp12_v_b_20')
// (30, 23, 'sp4_h_l_38')
// (30, 23, 'sp4_v_b_10')
// (30, 24, 'sp12_v_b_19')
// (30, 25, 'sp12_v_b_16')
// (30, 25, 'sp4_h_l_45')
// (30, 25, 'sp4_v_t_45')
// (30, 26, 'sp12_v_b_15')
// (30, 26, 'sp4_v_b_45')
// (30, 27, 'sp12_v_b_12')
// (30, 27, 'sp4_v_b_32')
// (30, 28, 'sp12_v_b_11')
// (30, 28, 'sp4_v_b_21')
// (30, 29, 'sp12_h_l_23')
// (30, 29, 'sp12_v_b_8')
// (30, 29, 'sp12_v_t_23')
// (30, 29, 'sp4_h_l_45')
// (30, 29, 'sp4_v_b_8')
// (30, 29, 'sp4_v_t_45')
// (30, 30, 'sp12_v_b_23')
// (30, 30, 'sp12_v_b_7')
// (30, 30, 'sp4_v_b_45')
// (30, 31, 'sp12_v_b_20')
// (30, 31, 'sp12_v_b_4')
// (30, 31, 'sp4_v_b_32')
// (30, 32, 'neigh_op_top_0')
// (30, 32, 'neigh_op_top_4')
// (30, 32, 'sp12_v_b_19')
// (30, 32, 'sp12_v_b_3')
// (30, 32, 'sp4_v_b_21')
// (30, 33, 'io_0/D_IN_0')
// (30, 33, 'io_0/PAD')
// (30, 33, 'span12_vert_0')
// (30, 33, 'span12_vert_16')
// (30, 33, 'span4_vert_8')
// (31, 32, 'neigh_op_tnl_0')
// (31, 32, 'neigh_op_tnl_4')

wire n48;
// (6, 22, 'neigh_op_tnr_5')
// (6, 23, 'neigh_op_rgt_5')
// (6, 24, 'neigh_op_bnr_5')
// (7, 22, 'neigh_op_top_5')
// (7, 23, 'local_g0_5')
// (7, 23, 'lutff_5/out')
// (7, 23, 'lutff_6/in_3')
// (7, 24, 'neigh_op_bot_5')
// (8, 22, 'neigh_op_tnl_5')
// (8, 23, 'neigh_op_lft_5')
// (8, 24, 'neigh_op_bnl_5')

wire n49;
// (6, 22, 'neigh_op_tnr_6')
// (6, 23, 'neigh_op_rgt_6')
// (6, 24, 'neigh_op_bnr_6')
// (7, 22, 'local_g1_6')
// (7, 22, 'lutff_1/in_0')
// (7, 22, 'neigh_op_top_6')
// (7, 23, 'lutff_6/out')
// (7, 24, 'neigh_op_bot_6')
// (8, 22, 'neigh_op_tnl_6')
// (8, 23, 'neigh_op_lft_6')
// (8, 24, 'neigh_op_bnl_6')

wire n50;
// (6, 22, 'sp4_r_v_b_37')
// (6, 23, 'sp4_r_v_b_24')
// (6, 24, 'neigh_op_tnr_0')
// (6, 24, 'sp4_r_v_b_13')
// (6, 25, 'neigh_op_rgt_0')
// (6, 25, 'sp4_r_v_b_0')
// (6, 26, 'neigh_op_bnr_0')
// (7, 21, 'local_g1_5')
// (7, 21, 'lutff_4/in_0')
// (7, 21, 'sp4_h_r_5')
// (7, 21, 'sp4_v_t_37')
// (7, 22, 'sp4_v_b_37')
// (7, 23, 'sp4_v_b_24')
// (7, 24, 'neigh_op_top_0')
// (7, 24, 'sp4_v_b_13')
// (7, 25, 'lutff_0/out')
// (7, 25, 'sp4_v_b_0')
// (7, 26, 'neigh_op_bot_0')
// (8, 21, 'sp4_h_r_16')
// (8, 24, 'neigh_op_tnl_0')
// (8, 25, 'neigh_op_lft_0')
// (8, 26, 'neigh_op_bnl_0')
// (9, 21, 'sp4_h_r_29')
// (10, 21, 'sp4_h_r_40')
// (11, 21, 'sp4_h_l_40')

wire io_33_30_0;
// (7, 13, 'sp4_r_v_b_38')
// (7, 14, 'sp4_r_v_b_27')
// (7, 15, 'sp4_r_v_b_14')
// (7, 15, 'sp4_r_v_b_36')
// (7, 16, 'sp4_r_v_b_25')
// (7, 16, 'sp4_r_v_b_3')
// (7, 17, 'sp4_r_v_b_12')
// (7, 17, 'sp4_r_v_b_41')
// (7, 18, 'sp4_r_v_b_1')
// (7, 18, 'sp4_r_v_b_28')
// (7, 19, 'sp4_r_v_b_17')
// (7, 19, 'sp4_r_v_b_39')
// (7, 20, 'sp4_r_v_b_26')
// (7, 20, 'sp4_r_v_b_4')
// (7, 21, 'sp4_r_v_b_15')
// (7, 21, 'sp4_r_v_b_47')
// (7, 22, 'sp4_r_v_b_2')
// (7, 22, 'sp4_r_v_b_34')
// (7, 23, 'sp4_r_v_b_23')
// (7, 23, 'sp4_r_v_b_42')
// (7, 24, 'sp4_r_v_b_10')
// (7, 24, 'sp4_r_v_b_31')
// (7, 25, 'sp4_r_v_b_18')
// (7, 26, 'sp4_r_v_b_7')
// (8, 12, 'sp4_v_t_38')
// (8, 13, 'sp4_v_b_38')
// (8, 14, 'sp4_v_b_27')
// (8, 14, 'sp4_v_t_36')
// (8, 15, 'local_g0_6')
// (8, 15, 'ram/RADDR_9')
// (8, 15, 'sp4_v_b_14')
// (8, 15, 'sp4_v_b_36')
// (8, 16, 'sp4_h_r_10')
// (8, 16, 'sp4_v_b_25')
// (8, 16, 'sp4_v_b_3')
// (8, 16, 'sp4_v_t_41')
// (8, 17, 'local_g0_4')
// (8, 17, 'ram/RADDR_9')
// (8, 17, 'sp4_v_b_12')
// (8, 17, 'sp4_v_b_41')
// (8, 18, 'sp12_v_t_23')
// (8, 18, 'sp4_h_r_8')
// (8, 18, 'sp4_v_b_1')
// (8, 18, 'sp4_v_b_28')
// (8, 18, 'sp4_v_t_39')
// (8, 19, 'local_g1_1')
// (8, 19, 'ram/RADDR_9')
// (8, 19, 'sp12_v_b_23')
// (8, 19, 'sp4_v_b_17')
// (8, 19, 'sp4_v_b_39')
// (8, 20, 'sp12_v_b_20')
// (8, 20, 'sp4_h_r_10')
// (8, 20, 'sp4_v_b_26')
// (8, 20, 'sp4_v_b_4')
// (8, 20, 'sp4_v_t_47')
// (8, 21, 'local_g1_7')
// (8, 21, 'ram/RADDR_9')
// (8, 21, 'sp12_v_b_19')
// (8, 21, 'sp4_v_b_15')
// (8, 21, 'sp4_v_b_47')
// (8, 22, 'sp12_v_b_16')
// (8, 22, 'sp4_h_r_1')
// (8, 22, 'sp4_v_b_2')
// (8, 22, 'sp4_v_b_34')
// (8, 22, 'sp4_v_t_42')
// (8, 23, 'local_g1_7')
// (8, 23, 'ram/RADDR_9')
// (8, 23, 'sp12_v_b_15')
// (8, 23, 'sp4_v_b_23')
// (8, 23, 'sp4_v_b_42')
// (8, 24, 'sp12_v_b_12')
// (8, 24, 'sp4_v_b_10')
// (8, 24, 'sp4_v_b_31')
// (8, 25, 'local_g0_2')
// (8, 25, 'ram/RADDR_9')
// (8, 25, 'sp12_v_b_11')
// (8, 25, 'sp4_v_b_18')
// (8, 26, 'sp12_v_b_8')
// (8, 26, 'sp4_v_b_7')
// (8, 27, 'local_g3_7')
// (8, 27, 'ram/RADDR_9')
// (8, 27, 'sp12_v_b_7')
// (8, 27, 'sp4_r_v_b_41')
// (8, 28, 'sp12_v_b_4')
// (8, 28, 'sp4_r_v_b_28')
// (8, 29, 'local_g3_1')
// (8, 29, 'ram/RADDR_9')
// (8, 29, 'sp12_v_b_3')
// (8, 29, 'sp4_r_v_b_17')
// (8, 30, 'sp12_h_r_0')
// (8, 30, 'sp12_v_b_0')
// (8, 30, 'sp4_r_v_b_4')
// (9, 16, 'sp4_h_r_23')
// (9, 18, 'sp4_h_r_21')
// (9, 20, 'sp4_h_r_23')
// (9, 22, 'sp4_h_r_12')
// (9, 26, 'sp4_v_t_41')
// (9, 27, 'sp4_v_b_41')
// (9, 28, 'sp4_v_b_28')
// (9, 29, 'sp4_v_b_17')
// (9, 30, 'sp12_h_r_3')
// (9, 30, 'sp4_h_r_11')
// (9, 30, 'sp4_v_b_4')
// (10, 16, 'sp4_h_r_34')
// (10, 18, 'sp4_h_r_32')
// (10, 20, 'sp4_h_r_34')
// (10, 22, 'sp4_h_r_25')
// (10, 30, 'sp12_h_r_4')
// (10, 30, 'sp4_h_r_22')
// (11, 16, 'sp4_h_r_47')
// (11, 17, 'sp4_r_v_b_47')
// (11, 18, 'sp4_h_r_45')
// (11, 18, 'sp4_r_v_b_34')
// (11, 19, 'sp4_r_v_b_23')
// (11, 19, 'sp4_r_v_b_45')
// (11, 20, 'sp4_h_r_47')
// (11, 20, 'sp4_r_v_b_10')
// (11, 20, 'sp4_r_v_b_32')
// (11, 21, 'sp4_r_v_b_21')
// (11, 22, 'sp4_h_r_36')
// (11, 22, 'sp4_r_v_b_8')
// (11, 30, 'sp12_h_r_7')
// (11, 30, 'sp4_h_r_35')
// (12, 16, 'sp4_h_l_47')
// (12, 16, 'sp4_v_t_47')
// (12, 17, 'sp4_v_b_47')
// (12, 18, 'sp12_v_t_23')
// (12, 18, 'sp4_h_l_45')
// (12, 18, 'sp4_v_b_34')
// (12, 18, 'sp4_v_t_45')
// (12, 19, 'sp12_v_b_23')
// (12, 19, 'sp4_v_b_23')
// (12, 19, 'sp4_v_b_45')
// (12, 20, 'sp12_v_b_20')
// (12, 20, 'sp4_h_l_47')
// (12, 20, 'sp4_v_b_10')
// (12, 20, 'sp4_v_b_32')
// (12, 21, 'sp12_v_b_19')
// (12, 21, 'sp4_v_b_21')
// (12, 22, 'sp12_v_b_16')
// (12, 22, 'sp4_h_l_36')
// (12, 22, 'sp4_v_b_8')
// (12, 23, 'sp12_v_b_15')
// (12, 24, 'sp12_v_b_12')
// (12, 25, 'sp12_v_b_11')
// (12, 26, 'sp12_v_b_8')
// (12, 27, 'sp12_v_b_7')
// (12, 28, 'sp12_v_b_4')
// (12, 29, 'sp12_v_b_3')
// (12, 30, 'sp12_h_r_0')
// (12, 30, 'sp12_h_r_8')
// (12, 30, 'sp12_v_b_0')
// (12, 30, 'sp4_h_r_46')
// (13, 30, 'sp12_h_r_11')
// (13, 30, 'sp12_h_r_3')
// (13, 30, 'sp4_h_l_46')
// (13, 30, 'sp4_h_r_3')
// (14, 30, 'sp12_h_r_12')
// (14, 30, 'sp12_h_r_4')
// (14, 30, 'sp4_h_r_14')
// (15, 30, 'sp12_h_r_15')
// (15, 30, 'sp12_h_r_7')
// (15, 30, 'sp4_h_r_27')
// (16, 30, 'sp12_h_r_16')
// (16, 30, 'sp12_h_r_8')
// (16, 30, 'sp4_h_r_38')
// (17, 30, 'sp12_h_r_11')
// (17, 30, 'sp12_h_r_19')
// (17, 30, 'sp4_h_l_38')
// (18, 30, 'sp12_h_r_12')
// (18, 30, 'sp12_h_r_20')
// (19, 30, 'sp12_h_r_15')
// (19, 30, 'sp12_h_r_23')
// (20, 20, 'local_g0_3')
// (20, 20, 'lutff_2/in_3')
// (20, 20, 'sp4_h_r_3')
// (20, 30, 'sp12_h_l_23')
// (20, 30, 'sp12_h_r_0')
// (20, 30, 'sp12_h_r_16')
// (21, 20, 'sp4_h_r_14')
// (21, 30, 'sp12_h_r_19')
// (21, 30, 'sp12_h_r_3')
// (22, 20, 'sp4_h_r_27')
// (22, 30, 'sp12_h_r_20')
// (22, 30, 'sp12_h_r_4')
// (23, 17, 'sp4_r_v_b_47')
// (23, 18, 'sp4_r_v_b_34')
// (23, 19, 'sp4_r_v_b_23')
// (23, 20, 'sp4_h_r_38')
// (23, 20, 'sp4_r_v_b_10')
// (23, 30, 'sp12_h_r_23')
// (23, 30, 'sp12_h_r_7')
// (24, 16, 'sp4_v_t_47')
// (24, 17, 'sp4_v_b_47')
// (24, 18, 'sp12_v_t_23')
// (24, 18, 'sp4_v_b_34')
// (24, 19, 'sp12_v_b_23')
// (24, 19, 'sp4_v_b_23')
// (24, 20, 'sp12_v_b_20')
// (24, 20, 'sp4_h_l_38')
// (24, 20, 'sp4_v_b_10')
// (24, 21, 'sp12_v_b_19')
// (24, 22, 'sp12_v_b_16')
// (24, 23, 'sp12_v_b_15')
// (24, 24, 'sp12_v_b_12')
// (24, 25, 'sp12_v_b_11')
// (24, 26, 'sp12_v_b_8')
// (24, 27, 'sp12_v_b_7')
// (24, 27, 'sp4_r_v_b_36')
// (24, 27, 'sp4_r_v_b_47')
// (24, 28, 'sp12_v_b_4')
// (24, 28, 'sp4_r_v_b_25')
// (24, 28, 'sp4_r_v_b_34')
// (24, 29, 'sp12_v_b_3')
// (24, 29, 'sp4_r_v_b_12')
// (24, 29, 'sp4_r_v_b_23')
// (24, 30, 'sp12_h_l_23')
// (24, 30, 'sp12_h_r_0')
// (24, 30, 'sp12_h_r_8')
// (24, 30, 'sp12_v_b_0')
// (24, 30, 'sp4_r_v_b_1')
// (24, 30, 'sp4_r_v_b_10')
// (25, 15, 'local_g3_3')
// (25, 15, 'ram/RADDR_9')
// (25, 15, 'sp4_r_v_b_43')
// (25, 16, 'sp4_r_v_b_30')
// (25, 17, 'local_g3_3')
// (25, 17, 'ram/RADDR_9')
// (25, 17, 'sp4_r_v_b_19')
// (25, 18, 'sp4_r_v_b_6')
// (25, 19, 'local_g3_3')
// (25, 19, 'ram/RADDR_9')
// (25, 19, 'sp4_r_v_b_43')
// (25, 20, 'sp4_r_v_b_30')
// (25, 21, 'local_g3_3')
// (25, 21, 'ram/RADDR_9')
// (25, 21, 'sp4_r_v_b_19')
// (25, 22, 'sp4_r_v_b_6')
// (25, 23, 'local_g2_4')
// (25, 23, 'ram/RADDR_9')
// (25, 23, 'sp4_r_v_b_36')
// (25, 24, 'sp4_r_v_b_25')
// (25, 25, 'local_g2_4')
// (25, 25, 'ram/RADDR_9')
// (25, 25, 'sp4_r_v_b_12')
// (25, 26, 'sp4_r_v_b_1')
// (25, 26, 'sp4_v_t_36')
// (25, 26, 'sp4_v_t_47')
// (25, 27, 'local_g2_4')
// (25, 27, 'ram/RADDR_9')
// (25, 27, 'sp4_v_b_36')
// (25, 27, 'sp4_v_b_47')
// (25, 28, 'sp4_v_b_25')
// (25, 28, 'sp4_v_b_34')
// (25, 29, 'local_g1_7')
// (25, 29, 'ram/RADDR_9')
// (25, 29, 'sp4_v_b_12')
// (25, 29, 'sp4_v_b_23')
// (25, 30, 'sp12_h_r_11')
// (25, 30, 'sp12_h_r_3')
// (25, 30, 'sp4_h_r_5')
// (25, 30, 'sp4_h_r_8')
// (25, 30, 'sp4_v_b_1')
// (25, 30, 'sp4_v_b_10')
// (26, 14, 'sp4_v_t_43')
// (26, 15, 'sp4_v_b_43')
// (26, 16, 'sp4_v_b_30')
// (26, 17, 'sp4_v_b_19')
// (26, 18, 'sp4_h_r_1')
// (26, 18, 'sp4_v_b_6')
// (26, 18, 'sp4_v_t_43')
// (26, 19, 'sp4_v_b_43')
// (26, 20, 'sp4_v_b_30')
// (26, 21, 'local_g0_3')
// (26, 21, 'lutff_2/in_3')
// (26, 21, 'sp4_v_b_19')
// (26, 22, 'sp4_h_r_1')
// (26, 22, 'sp4_v_b_6')
// (26, 22, 'sp4_v_t_36')
// (26, 23, 'sp4_v_b_36')
// (26, 24, 'sp4_v_b_25')
// (26, 25, 'sp4_v_b_12')
// (26, 26, 'sp4_h_r_1')
// (26, 26, 'sp4_v_b_1')
// (26, 30, 'sp12_h_r_12')
// (26, 30, 'sp12_h_r_4')
// (26, 30, 'sp4_h_r_16')
// (26, 30, 'sp4_h_r_21')
// (27, 18, 'sp4_h_r_12')
// (27, 22, 'sp4_h_r_12')
// (27, 26, 'sp4_h_r_12')
// (27, 30, 'sp12_h_r_15')
// (27, 30, 'sp12_h_r_7')
// (27, 30, 'sp4_h_r_29')
// (27, 30, 'sp4_h_r_32')
// (28, 18, 'sp4_h_r_25')
// (28, 22, 'sp4_h_r_25')
// (28, 26, 'sp4_h_r_25')
// (28, 30, 'sp12_h_r_16')
// (28, 30, 'sp12_h_r_8')
// (28, 30, 'sp4_h_r_40')
// (28, 30, 'sp4_h_r_45')
// (29, 18, 'sp4_h_r_36')
// (29, 22, 'sp4_h_r_36')
// (29, 26, 'sp4_h_r_36')
// (29, 30, 'sp12_h_r_11')
// (29, 30, 'sp12_h_r_19')
// (29, 30, 'sp4_h_l_40')
// (29, 30, 'sp4_h_l_45')
// (29, 30, 'sp4_h_r_5')
// (30, 18, 'sp4_h_l_36')
// (30, 18, 'sp4_h_r_1')
// (30, 22, 'sp4_h_l_36')
// (30, 22, 'sp4_h_r_1')
// (30, 26, 'sp4_h_l_36')
// (30, 26, 'sp4_h_r_1')
// (30, 30, 'sp12_h_r_12')
// (30, 30, 'sp12_h_r_20')
// (30, 30, 'sp4_h_r_16')
// (31, 18, 'sp4_h_r_12')
// (31, 22, 'sp4_h_r_12')
// (31, 26, 'sp4_h_r_12')
// (31, 30, 'sp12_h_r_15')
// (31, 30, 'sp12_h_r_23')
// (31, 30, 'sp4_h_r_29')
// (32, 18, 'sp4_h_r_25')
// (32, 22, 'sp4_h_r_25')
// (32, 26, 'sp4_h_r_25')
// (32, 29, 'neigh_op_tnr_0')
// (32, 29, 'neigh_op_tnr_4')
// (32, 30, 'neigh_op_rgt_0')
// (32, 30, 'neigh_op_rgt_4')
// (32, 30, 'sp12_h_l_23')
// (32, 30, 'sp12_h_r_0')
// (32, 30, 'sp12_h_r_16')
// (32, 30, 'sp4_h_r_40')
// (32, 31, 'neigh_op_bnr_0')
// (32, 31, 'neigh_op_bnr_4')
// (33, 18, 'span4_horz_25')
// (33, 18, 'span4_vert_t_12')
// (33, 19, 'span4_vert_b_12')
// (33, 20, 'span4_vert_b_8')
// (33, 21, 'span4_vert_b_4')
// (33, 22, 'span4_horz_25')
// (33, 22, 'span4_vert_b_0')
// (33, 22, 'span4_vert_t_12')
// (33, 23, 'span4_vert_b_12')
// (33, 24, 'span4_vert_b_8')
// (33, 25, 'span4_vert_b_4')
// (33, 26, 'span4_horz_25')
// (33, 26, 'span4_vert_b_0')
// (33, 26, 'span4_vert_t_12')
// (33, 27, 'span4_vert_b_12')
// (33, 28, 'span4_vert_b_8')
// (33, 29, 'span4_vert_b_4')
// (33, 30, 'io_0/D_IN_0')
// (33, 30, 'io_0/PAD')
// (33, 30, 'span12_horz_0')
// (33, 30, 'span12_horz_16')
// (33, 30, 'span4_horz_40')
// (33, 30, 'span4_vert_b_0')

wire n52;
// (7, 13, 'sp4_r_v_b_42')
// (7, 14, 'sp4_r_v_b_31')
// (7, 15, 'sp4_r_v_b_18')
// (7, 16, 'sp4_r_v_b_7')
// (8, 12, 'sp4_v_t_42')
// (8, 13, 'sp4_v_b_42')
// (8, 14, 'sp4_v_b_31')
// (8, 15, 'local_g0_2')
// (8, 15, 'ram/RCLKE')
// (8, 15, 'sp4_v_b_18')
// (8, 16, 'sp4_h_r_7')
// (8, 16, 'sp4_v_b_7')
// (9, 16, 'sp4_h_r_18')
// (10, 16, 'sp4_h_r_31')
// (11, 16, 'sp4_h_r_42')
// (12, 16, 'sp4_h_l_42')
// (12, 16, 'sp4_h_r_11')
// (13, 16, 'sp4_h_r_22')
// (14, 16, 'sp4_h_r_35')
// (15, 16, 'sp4_h_r_46')
// (16, 16, 'sp4_h_l_46')
// (16, 16, 'sp4_h_r_11')
// (17, 16, 'sp4_h_r_22')
// (17, 21, 'sp4_r_v_b_41')
// (17, 22, 'sp4_r_v_b_28')
// (17, 23, 'sp4_r_v_b_17')
// (17, 24, 'sp4_r_v_b_4')
// (18, 16, 'sp4_h_r_35')
// (18, 20, 'sp4_h_r_10')
// (18, 20, 'sp4_v_t_41')
// (18, 21, 'sp4_v_b_41')
// (18, 22, 'sp4_v_b_28')
// (18, 23, 'local_g0_1')
// (18, 23, 'lutff_7/in_2')
// (18, 23, 'sp4_v_b_17')
// (18, 24, 'sp4_v_b_4')
// (19, 16, 'sp4_h_r_46')
// (19, 20, 'sp4_h_r_23')
// (20, 16, 'sp4_h_l_46')
// (20, 16, 'sp4_h_r_8')
// (20, 20, 'sp4_h_r_34')
// (21, 16, 'sp4_h_r_21')
// (21, 20, 'sp4_h_r_47')
// (22, 16, 'sp4_h_r_32')
// (22, 20, 'sp4_h_l_47')
// (22, 20, 'sp4_h_r_10')
// (23, 16, 'sp4_h_r_45')
// (23, 17, 'sp4_r_v_b_39')
// (23, 18, 'sp4_r_v_b_26')
// (23, 18, 'sp4_r_v_b_42')
// (23, 19, 'neigh_op_tnr_1')
// (23, 19, 'sp4_r_v_b_15')
// (23, 19, 'sp4_r_v_b_31')
// (23, 20, 'neigh_op_rgt_1')
// (23, 20, 'sp4_h_r_23')
// (23, 20, 'sp4_r_v_b_18')
// (23, 20, 'sp4_r_v_b_2')
// (23, 21, 'neigh_op_bnr_1')
// (23, 21, 'sp4_r_v_b_7')
// (24, 13, 'sp4_r_v_b_43')
// (24, 14, 'sp4_r_v_b_30')
// (24, 15, 'sp4_r_v_b_19')
// (24, 16, 'sp4_h_l_45')
// (24, 16, 'sp4_r_v_b_6')
// (24, 16, 'sp4_v_t_39')
// (24, 17, 'sp4_r_v_b_38')
// (24, 17, 'sp4_v_b_39')
// (24, 17, 'sp4_v_t_42')
// (24, 18, 'sp4_r_v_b_27')
// (24, 18, 'sp4_v_b_26')
// (24, 18, 'sp4_v_b_42')
// (24, 19, 'neigh_op_top_1')
// (24, 19, 'sp4_r_v_b_14')
// (24, 19, 'sp4_r_v_b_46')
// (24, 19, 'sp4_v_b_15')
// (24, 19, 'sp4_v_b_31')
// (24, 20, 'lutff_1/out')
// (24, 20, 'sp4_h_r_34')
// (24, 20, 'sp4_r_v_b_3')
// (24, 20, 'sp4_r_v_b_35')
// (24, 20, 'sp4_v_b_18')
// (24, 20, 'sp4_v_b_2')
// (24, 21, 'neigh_op_bot_1')
// (24, 21, 'sp4_h_r_7')
// (24, 21, 'sp4_r_v_b_22')
// (24, 21, 'sp4_v_b_7')
// (24, 22, 'sp4_r_v_b_11')
// (24, 23, 'sp4_r_v_b_42')
// (24, 24, 'sp4_r_v_b_31')
// (24, 25, 'sp4_r_v_b_18')
// (24, 26, 'sp4_r_v_b_7')
// (25, 12, 'sp4_v_t_43')
// (25, 13, 'sp4_v_b_43')
// (25, 14, 'sp4_v_b_30')
// (25, 15, 'local_g1_3')
// (25, 15, 'ram/RCLKE')
// (25, 15, 'sp4_v_b_19')
// (25, 16, 'sp4_v_b_6')
// (25, 16, 'sp4_v_t_38')
// (25, 17, 'sp4_v_b_38')
// (25, 18, 'sp4_v_b_27')
// (25, 18, 'sp4_v_t_46')
// (25, 19, 'neigh_op_tnl_1')
// (25, 19, 'sp4_v_b_14')
// (25, 19, 'sp4_v_b_46')
// (25, 20, 'neigh_op_lft_1')
// (25, 20, 'sp4_h_r_47')
// (25, 20, 'sp4_v_b_3')
// (25, 20, 'sp4_v_b_35')
// (25, 21, 'local_g0_2')
// (25, 21, 'neigh_op_bnl_1')
// (25, 21, 'ram/RCLKE')
// (25, 21, 'sp4_h_r_18')
// (25, 21, 'sp4_v_b_22')
// (25, 22, 'sp4_v_b_11')
// (25, 22, 'sp4_v_t_42')
// (25, 23, 'sp4_v_b_42')
// (25, 24, 'sp4_v_b_31')
// (25, 25, 'local_g0_2')
// (25, 25, 'ram/RCLKE')
// (25, 25, 'sp4_v_b_18')
// (25, 26, 'sp4_v_b_7')
// (26, 20, 'sp4_h_l_47')
// (26, 21, 'sp4_h_r_31')
// (27, 21, 'sp4_h_r_42')
// (28, 21, 'sp4_h_l_42')

wire n53;
// (7, 14, 'neigh_op_tnr_4')
// (7, 15, 'neigh_op_rgt_4')
// (7, 16, 'neigh_op_bnr_4')
// (8, 12, 'sp4_r_v_b_44')
// (8, 13, 'sp4_r_v_b_33')
// (8, 14, 'neigh_op_top_4')
// (8, 14, 'sp4_r_v_b_20')
// (8, 15, 'ram/RDATA_11')
// (8, 15, 'sp4_r_v_b_9')
// (8, 16, 'neigh_op_bot_4')
// (8, 16, 'sp4_r_v_b_40')
// (8, 17, 'sp4_r_v_b_29')
// (8, 18, 'sp4_r_v_b_16')
// (8, 19, 'sp4_r_v_b_5')
// (9, 11, 'sp4_v_t_44')
// (9, 12, 'sp4_v_b_44')
// (9, 13, 'sp4_v_b_33')
// (9, 14, 'neigh_op_tnl_4')
// (9, 14, 'sp4_v_b_20')
// (9, 15, 'neigh_op_lft_4')
// (9, 15, 'sp4_v_b_9')
// (9, 15, 'sp4_v_t_40')
// (9, 16, 'neigh_op_bnl_4')
// (9, 16, 'sp4_v_b_40')
// (9, 17, 'sp4_v_b_29')
// (9, 18, 'sp4_v_b_16')
// (9, 19, 'local_g0_5')
// (9, 19, 'lutff_0/in_1')
// (9, 19, 'sp4_v_b_5')

wire n54;
// (7, 15, 'neigh_op_tnr_4')
// (7, 16, 'neigh_op_rgt_4')
// (7, 17, 'neigh_op_bnr_4')
// (8, 15, 'neigh_op_top_4')
// (8, 16, 'ram/RDATA_3')
// (8, 16, 'sp4_r_v_b_41')
// (8, 17, 'neigh_op_bot_4')
// (8, 17, 'sp4_r_v_b_28')
// (8, 18, 'sp4_r_v_b_17')
// (8, 19, 'sp4_r_v_b_4')
// (9, 15, 'neigh_op_tnl_4')
// (9, 15, 'sp4_v_t_41')
// (9, 16, 'neigh_op_lft_4')
// (9, 16, 'sp4_v_b_41')
// (9, 17, 'neigh_op_bnl_4')
// (9, 17, 'sp4_v_b_28')
// (9, 18, 'sp4_v_b_17')
// (9, 19, 'local_g1_4')
// (9, 19, 'lutff_1/in_2')
// (9, 19, 'sp4_v_b_4')

wire io_33_27_1;
// (7, 15, 'sp4_h_r_3')
// (7, 19, 'sp4_h_r_3')
// (7, 27, 'sp4_h_r_11')
// (8, 15, 'local_g1_6')
// (8, 15, 'ram/RADDR_10')
// (8, 15, 'sp4_h_r_14')
// (8, 16, 'sp4_r_v_b_42')
// (8, 17, 'local_g0_7')
// (8, 17, 'ram/RADDR_10')
// (8, 17, 'sp4_r_v_b_31')
// (8, 18, 'sp4_r_v_b_18')
// (8, 19, 'local_g1_6')
// (8, 19, 'ram/RADDR_10')
// (8, 19, 'sp4_h_r_14')
// (8, 19, 'sp4_r_v_b_7')
// (8, 20, 'sp4_r_v_b_41')
// (8, 20, 'sp4_r_v_b_44')
// (8, 21, 'local_g1_4')
// (8, 21, 'ram/RADDR_10')
// (8, 21, 'sp4_r_v_b_28')
// (8, 21, 'sp4_r_v_b_33')
// (8, 22, 'sp4_r_v_b_17')
// (8, 22, 'sp4_r_v_b_20')
// (8, 23, 'local_g2_1')
// (8, 23, 'ram/RADDR_10')
// (8, 23, 'sp4_r_v_b_4')
// (8, 23, 'sp4_r_v_b_9')
// (8, 24, 'sp4_r_v_b_36')
// (8, 25, 'local_g0_1')
// (8, 25, 'ram/RADDR_10')
// (8, 25, 'sp4_r_v_b_25')
// (8, 26, 'sp4_r_v_b_12')
// (8, 27, 'local_g1_6')
// (8, 27, 'ram/RADDR_10')
// (8, 27, 'sp4_h_r_22')
// (8, 27, 'sp4_r_v_b_1')
// (8, 28, 'sp4_r_v_b_36')
// (8, 29, 'local_g0_1')
// (8, 29, 'ram/RADDR_10')
// (8, 29, 'sp4_r_v_b_25')
// (8, 30, 'sp4_r_v_b_12')
// (8, 31, 'sp4_r_v_b_1')
// (9, 15, 'sp4_h_r_1')
// (9, 15, 'sp4_h_r_27')
// (9, 15, 'sp4_v_t_42')
// (9, 16, 'sp4_v_b_42')
// (9, 17, 'sp4_v_b_31')
// (9, 18, 'sp4_v_b_18')
// (9, 19, 'sp4_h_r_27')
// (9, 19, 'sp4_v_b_7')
// (9, 19, 'sp4_v_t_41')
// (9, 19, 'sp4_v_t_44')
// (9, 20, 'sp4_v_b_41')
// (9, 20, 'sp4_v_b_44')
// (9, 21, 'sp4_v_b_28')
// (9, 21, 'sp4_v_b_33')
// (9, 22, 'sp4_v_b_17')
// (9, 22, 'sp4_v_b_20')
// (9, 23, 'sp4_v_b_4')
// (9, 23, 'sp4_v_b_9')
// (9, 23, 'sp4_v_t_36')
// (9, 24, 'sp4_v_b_36')
// (9, 25, 'sp4_v_b_25')
// (9, 26, 'sp4_v_b_12')
// (9, 27, 'sp4_h_r_1')
// (9, 27, 'sp4_h_r_35')
// (9, 27, 'sp4_v_b_1')
// (9, 27, 'sp4_v_t_36')
// (9, 28, 'sp4_v_b_36')
// (9, 29, 'sp4_v_b_25')
// (9, 30, 'sp4_v_b_12')
// (9, 31, 'sp4_v_b_1')
// (10, 15, 'sp12_h_r_0')
// (10, 15, 'sp4_h_r_12')
// (10, 15, 'sp4_h_r_38')
// (10, 16, 'sp4_r_v_b_38')
// (10, 17, 'sp4_r_v_b_27')
// (10, 18, 'sp4_r_v_b_14')
// (10, 19, 'sp4_h_r_38')
// (10, 19, 'sp4_r_v_b_3')
// (10, 27, 'sp12_h_r_0')
// (10, 27, 'sp4_h_r_12')
// (10, 27, 'sp4_h_r_46')
// (11, 15, 'sp12_h_r_3')
// (11, 15, 'sp4_h_l_38')
// (11, 15, 'sp4_h_r_25')
// (11, 15, 'sp4_h_r_3')
// (11, 15, 'sp4_v_t_38')
// (11, 16, 'sp4_v_b_38')
// (11, 17, 'sp4_v_b_27')
// (11, 18, 'sp4_v_b_14')
// (11, 19, 'sp4_h_l_38')
// (11, 19, 'sp4_v_b_3')
// (11, 27, 'sp12_h_r_3')
// (11, 27, 'sp4_h_l_46')
// (11, 27, 'sp4_h_r_25')
// (11, 27, 'sp4_h_r_3')
// (12, 15, 'sp12_h_r_4')
// (12, 15, 'sp4_h_r_14')
// (12, 15, 'sp4_h_r_36')
// (12, 27, 'sp12_h_r_4')
// (12, 27, 'sp4_h_r_14')
// (12, 27, 'sp4_h_r_36')
// (13, 15, 'sp12_h_r_7')
// (13, 15, 'sp4_h_l_36')
// (13, 15, 'sp4_h_r_27')
// (13, 27, 'sp12_h_r_7')
// (13, 27, 'sp4_h_l_36')
// (13, 27, 'sp4_h_r_27')
// (14, 15, 'sp12_h_r_8')
// (14, 15, 'sp4_h_r_38')
// (14, 27, 'sp12_h_r_8')
// (14, 27, 'sp4_h_r_38')
// (15, 15, 'sp12_h_r_11')
// (15, 15, 'sp4_h_l_38')
// (15, 27, 'sp12_h_r_11')
// (15, 27, 'sp4_h_l_38')
// (16, 15, 'sp12_h_r_12')
// (16, 27, 'sp12_h_r_12')
// (17, 15, 'sp12_h_r_15')
// (17, 27, 'sp12_h_r_15')
// (18, 15, 'sp12_h_r_16')
// (18, 27, 'sp12_h_r_16')
// (19, 15, 'sp12_h_r_19')
// (19, 27, 'sp12_h_r_19')
// (20, 15, 'sp12_h_r_20')
// (20, 27, 'sp12_h_r_20')
// (21, 15, 'sp12_h_r_23')
// (21, 27, 'sp12_h_r_23')
// (22, 15, 'sp12_h_l_23')
// (22, 15, 'sp12_v_t_23')
// (22, 16, 'sp12_v_b_23')
// (22, 17, 'sp12_v_b_20')
// (22, 18, 'sp12_v_b_19')
// (22, 19, 'sp12_v_b_16')
// (22, 20, 'sp12_v_b_15')
// (22, 21, 'local_g3_4')
// (22, 21, 'lutff_3/in_0')
// (22, 21, 'sp12_v_b_12')
// (22, 22, 'sp12_v_b_11')
// (22, 23, 'sp12_v_b_8')
// (22, 24, 'sp12_v_b_7')
// (22, 25, 'sp12_v_b_4')
// (22, 26, 'sp12_v_b_3')
// (22, 27, 'sp12_h_l_23')
// (22, 27, 'sp12_h_r_0')
// (22, 27, 'sp12_v_b_0')
// (23, 27, 'sp12_h_r_3')
// (24, 16, 'sp4_r_v_b_40')
// (24, 17, 'sp4_r_v_b_29')
// (24, 18, 'sp4_r_v_b_16')
// (24, 19, 'sp4_r_v_b_5')
// (24, 20, 'sp4_r_v_b_44')
// (24, 21, 'local_g2_1')
// (24, 21, 'lutff_2/in_1')
// (24, 21, 'sp4_r_v_b_33')
// (24, 22, 'sp4_r_v_b_20')
// (24, 23, 'sp4_r_v_b_9')
// (24, 24, 'sp4_r_v_b_40')
// (24, 25, 'sp4_r_v_b_29')
// (24, 26, 'sp4_r_v_b_16')
// (24, 27, 'sp12_h_r_4')
// (24, 27, 'sp4_r_v_b_5')
// (24, 28, 'sp4_r_v_b_43')
// (24, 29, 'sp4_r_v_b_30')
// (24, 30, 'sp4_r_v_b_19')
// (24, 31, 'sp4_r_v_b_6')
// (25, 15, 'local_g0_5')
// (25, 15, 'ram/RADDR_10')
// (25, 15, 'sp4_h_r_5')
// (25, 15, 'sp4_v_t_40')
// (25, 16, 'sp4_v_b_40')
// (25, 17, 'local_g2_5')
// (25, 17, 'ram/RADDR_10')
// (25, 17, 'sp4_v_b_29')
// (25, 18, 'sp4_v_b_16')
// (25, 19, 'local_g1_2')
// (25, 19, 'ram/RADDR_10')
// (25, 19, 'sp4_h_r_2')
// (25, 19, 'sp4_v_b_5')
// (25, 19, 'sp4_v_t_44')
// (25, 20, 'sp4_v_b_44')
// (25, 21, 'local_g2_1')
// (25, 21, 'ram/RADDR_10')
// (25, 21, 'sp4_v_b_33')
// (25, 22, 'sp4_v_b_20')
// (25, 23, 'local_g0_1')
// (25, 23, 'ram/RADDR_10')
// (25, 23, 'sp4_h_r_9')
// (25, 23, 'sp4_v_b_9')
// (25, 23, 'sp4_v_t_40')
// (25, 24, 'sp4_v_b_40')
// (25, 25, 'local_g2_5')
// (25, 25, 'ram/RADDR_10')
// (25, 25, 'sp4_v_b_29')
// (25, 26, 'sp4_v_b_16')
// (25, 27, 'local_g1_0')
// (25, 27, 'ram/RADDR_10')
// (25, 27, 'sp12_h_r_7')
// (25, 27, 'sp4_h_r_0')
// (25, 27, 'sp4_v_b_5')
// (25, 27, 'sp4_v_t_43')
// (25, 28, 'sp4_v_b_43')
// (25, 29, 'local_g3_6')
// (25, 29, 'ram/RADDR_10')
// (25, 29, 'sp4_v_b_30')
// (25, 30, 'sp4_v_b_19')
// (25, 31, 'sp4_v_b_6')
// (26, 15, 'sp4_h_r_16')
// (26, 19, 'sp4_h_r_15')
// (26, 23, 'sp4_h_r_20')
// (26, 27, 'sp12_h_r_8')
// (26, 27, 'sp4_h_r_13')
// (27, 15, 'sp4_h_r_29')
// (27, 19, 'sp4_h_r_26')
// (27, 23, 'sp4_h_r_33')
// (27, 27, 'sp12_h_r_11')
// (27, 27, 'sp4_h_r_24')
// (28, 15, 'sp4_h_r_40')
// (28, 19, 'sp4_h_r_39')
// (28, 23, 'sp4_h_r_44')
// (28, 24, 'sp4_r_v_b_44')
// (28, 25, 'sp4_r_v_b_33')
// (28, 26, 'sp4_r_v_b_20')
// (28, 27, 'sp12_h_r_12')
// (28, 27, 'sp4_h_r_37')
// (28, 27, 'sp4_r_v_b_9')
// (29, 15, 'sp4_h_l_40')
// (29, 19, 'sp4_h_l_39')
// (29, 23, 'sp4_h_l_44')
// (29, 23, 'sp4_v_t_44')
// (29, 24, 'sp4_v_b_44')
// (29, 25, 'sp4_v_b_33')
// (29, 26, 'sp4_v_b_20')
// (29, 27, 'sp12_h_r_15')
// (29, 27, 'sp4_h_l_37')
// (29, 27, 'sp4_h_r_9')
// (29, 27, 'sp4_v_b_9')
// (30, 27, 'sp12_h_r_16')
// (30, 27, 'sp4_h_r_20')
// (31, 27, 'sp12_h_r_19')
// (31, 27, 'sp4_h_r_33')
// (32, 26, 'neigh_op_tnr_2')
// (32, 26, 'neigh_op_tnr_6')
// (32, 27, 'neigh_op_rgt_2')
// (32, 27, 'neigh_op_rgt_6')
// (32, 27, 'sp12_h_r_20')
// (32, 27, 'sp4_h_r_44')
// (32, 28, 'neigh_op_bnr_2')
// (32, 28, 'neigh_op_bnr_6')
// (33, 27, 'io_1/D_IN_0')
// (33, 27, 'io_1/PAD')
// (33, 27, 'span12_horz_20')
// (33, 27, 'span4_horz_44')

wire n56;
// (7, 16, 'neigh_op_tnr_4')
// (7, 17, 'neigh_op_rgt_4')
// (7, 17, 'sp4_r_v_b_40')
// (7, 18, 'neigh_op_bnr_4')
// (7, 18, 'sp4_r_v_b_29')
// (7, 19, 'local_g3_0')
// (7, 19, 'lutff_2/in_3')
// (7, 19, 'sp4_r_v_b_16')
// (7, 20, 'sp4_r_v_b_5')
// (8, 16, 'neigh_op_top_4')
// (8, 16, 'sp4_v_t_40')
// (8, 17, 'ram/RDATA_11')
// (8, 17, 'sp4_v_b_40')
// (8, 18, 'neigh_op_bot_4')
// (8, 18, 'sp4_v_b_29')
// (8, 19, 'sp4_v_b_16')
// (8, 20, 'sp4_v_b_5')
// (9, 16, 'neigh_op_tnl_4')
// (9, 17, 'neigh_op_lft_4')
// (9, 18, 'neigh_op_bnl_4')

wire n57;
// (7, 17, 'neigh_op_tnr_4')
// (7, 18, 'neigh_op_rgt_4')
// (7, 19, 'local_g0_4')
// (7, 19, 'lutff_4/in_0')
// (7, 19, 'neigh_op_bnr_4')
// (8, 17, 'neigh_op_top_4')
// (8, 18, 'ram/RDATA_3')
// (8, 19, 'neigh_op_bot_4')
// (9, 17, 'neigh_op_tnl_4')
// (9, 18, 'neigh_op_lft_4')
// (9, 19, 'neigh_op_bnl_4')

reg n58 = 0;
// (7, 17, 'sp4_r_v_b_37')
// (7, 18, 'sp4_r_v_b_24')
// (7, 19, 'local_g2_5')
// (7, 19, 'lutff_2/in_1')
// (7, 19, 'sp4_r_v_b_13')
// (7, 20, 'sp4_r_v_b_0')
// (7, 21, 'sp4_r_v_b_37')
// (7, 21, 'sp4_r_v_b_43')
// (7, 22, 'sp4_r_v_b_24')
// (7, 22, 'sp4_r_v_b_30')
// (7, 23, 'local_g2_5')
// (7, 23, 'local_g3_3')
// (7, 23, 'lutff_0/in_2')
// (7, 23, 'lutff_5/in_0')
// (7, 23, 'sp4_r_v_b_13')
// (7, 23, 'sp4_r_v_b_19')
// (7, 23, 'sp4_r_v_b_37')
// (7, 24, 'sp4_r_v_b_0')
// (7, 24, 'sp4_r_v_b_24')
// (7, 24, 'sp4_r_v_b_6')
// (7, 25, 'local_g2_5')
// (7, 25, 'lutff_0/in_1')
// (7, 25, 'sp4_r_v_b_13')
// (7, 26, 'sp4_r_v_b_0')
// (8, 16, 'sp4_v_t_37')
// (8, 17, 'sp4_r_v_b_40')
// (8, 17, 'sp4_v_b_37')
// (8, 18, 'sp4_r_v_b_29')
// (8, 18, 'sp4_v_b_24')
// (8, 19, 'sp4_r_v_b_16')
// (8, 19, 'sp4_v_b_13')
// (8, 20, 'sp4_h_r_0')
// (8, 20, 'sp4_r_v_b_5')
// (8, 20, 'sp4_v_b_0')
// (8, 20, 'sp4_v_t_37')
// (8, 20, 'sp4_v_t_43')
// (8, 21, 'sp4_r_v_b_46')
// (8, 21, 'sp4_v_b_37')
// (8, 21, 'sp4_v_b_43')
// (8, 22, 'sp4_h_r_0')
// (8, 22, 'sp4_r_v_b_35')
// (8, 22, 'sp4_v_b_24')
// (8, 22, 'sp4_v_b_30')
// (8, 22, 'sp4_v_t_37')
// (8, 23, 'sp4_r_v_b_22')
// (8, 23, 'sp4_r_v_b_45')
// (8, 23, 'sp4_v_b_13')
// (8, 23, 'sp4_v_b_19')
// (8, 23, 'sp4_v_b_37')
// (8, 24, 'sp4_r_v_b_11')
// (8, 24, 'sp4_r_v_b_32')
// (8, 24, 'sp4_v_b_0')
// (8, 24, 'sp4_v_b_24')
// (8, 24, 'sp4_v_b_6')
// (8, 25, 'sp4_r_v_b_21')
// (8, 25, 'sp4_v_b_13')
// (8, 26, 'sp4_r_v_b_8')
// (8, 26, 'sp4_v_b_0')
// (9, 16, 'sp4_v_t_40')
// (9, 17, 'sp4_v_b_40')
// (9, 18, 'sp4_v_b_29')
// (9, 19, 'local_g1_0')
// (9, 19, 'lutff_2/in_1')
// (9, 19, 'sp4_v_b_16')
// (9, 20, 'sp4_h_r_13')
// (9, 20, 'sp4_h_r_5')
// (9, 20, 'sp4_v_b_5')
// (9, 20, 'sp4_v_t_46')
// (9, 21, 'sp4_v_b_46')
// (9, 22, 'sp4_h_r_13')
// (9, 22, 'sp4_h_r_2')
// (9, 22, 'sp4_v_b_35')
// (9, 22, 'sp4_v_t_45')
// (9, 23, 'local_g1_6')
// (9, 23, 'lutff_3/in_0')
// (9, 23, 'sp4_v_b_22')
// (9, 23, 'sp4_v_b_45')
// (9, 24, 'sp4_v_b_11')
// (9, 24, 'sp4_v_b_32')
// (9, 25, 'local_g0_5')
// (9, 25, 'lutff_6/in_1')
// (9, 25, 'sp4_v_b_21')
// (9, 26, 'sp4_v_b_8')
// (10, 20, 'sp4_h_r_16')
// (10, 20, 'sp4_h_r_24')
// (10, 22, 'sp4_h_r_15')
// (10, 22, 'sp4_h_r_24')
// (11, 20, 'sp4_h_r_29')
// (11, 20, 'sp4_h_r_37')
// (11, 22, 'sp4_h_r_26')
// (11, 22, 'sp4_h_r_37')
// (12, 20, 'sp4_h_l_37')
// (12, 20, 'sp4_h_r_4')
// (12, 20, 'sp4_h_r_40')
// (12, 22, 'sp4_h_l_37')
// (12, 22, 'sp4_h_r_0')
// (12, 22, 'sp4_h_r_39')
// (13, 20, 'sp4_h_l_40')
// (13, 20, 'sp4_h_r_17')
// (13, 20, 'sp4_h_r_5')
// (13, 22, 'sp4_h_l_39')
// (13, 22, 'sp4_h_r_13')
// (13, 22, 'sp4_h_r_6')
// (14, 20, 'sp4_h_r_16')
// (14, 20, 'sp4_h_r_28')
// (14, 22, 'sp4_h_r_19')
// (14, 22, 'sp4_h_r_24')
// (15, 19, 'neigh_op_tnr_4')
// (15, 19, 'sp4_r_v_b_37')
// (15, 20, 'neigh_op_rgt_4')
// (15, 20, 'sp4_h_r_29')
// (15, 20, 'sp4_h_r_41')
// (15, 20, 'sp4_r_v_b_24')
// (15, 21, 'neigh_op_bnr_4')
// (15, 21, 'sp4_r_v_b_13')
// (15, 22, 'sp4_h_r_30')
// (15, 22, 'sp4_h_r_37')
// (15, 22, 'sp4_r_v_b_0')
// (16, 18, 'sp4_v_t_37')
// (16, 19, 'neigh_op_top_4')
// (16, 19, 'sp4_r_v_b_36')
// (16, 19, 'sp4_v_b_37')
// (16, 20, 'lutff_4/out')
// (16, 20, 'sp4_h_l_41')
// (16, 20, 'sp4_h_r_40')
// (16, 20, 'sp4_h_r_8')
// (16, 20, 'sp4_r_v_b_25')
// (16, 20, 'sp4_r_v_b_41')
// (16, 20, 'sp4_v_b_24')
// (16, 21, 'neigh_op_bot_4')
// (16, 21, 'sp4_r_v_b_12')
// (16, 21, 'sp4_r_v_b_28')
// (16, 21, 'sp4_v_b_13')
// (16, 22, 'sp4_h_l_37')
// (16, 22, 'sp4_h_r_43')
// (16, 22, 'sp4_r_v_b_1')
// (16, 22, 'sp4_r_v_b_17')
// (16, 22, 'sp4_v_b_0')
// (16, 23, 'sp4_r_v_b_4')
// (17, 18, 'sp4_v_t_36')
// (17, 19, 'neigh_op_tnl_4')
// (17, 19, 'sp4_v_b_36')
// (17, 19, 'sp4_v_t_41')
// (17, 20, 'neigh_op_lft_4')
// (17, 20, 'sp4_h_l_40')
// (17, 20, 'sp4_h_r_21')
// (17, 20, 'sp4_v_b_25')
// (17, 20, 'sp4_v_b_41')
// (17, 21, 'neigh_op_bnl_4')
// (17, 21, 'sp4_v_b_12')
// (17, 21, 'sp4_v_b_28')
// (17, 22, 'sp4_h_l_43')
// (17, 22, 'sp4_v_b_1')
// (17, 22, 'sp4_v_b_17')
// (17, 23, 'sp4_h_r_10')
// (17, 23, 'sp4_v_b_4')
// (18, 20, 'sp4_h_r_32')
// (18, 23, 'sp4_h_r_23')
// (19, 20, 'sp4_h_r_45')
// (19, 23, 'sp4_h_r_34')
// (20, 20, 'sp4_h_l_45')
// (20, 23, 'sp4_h_r_47')
// (21, 23, 'sp4_h_l_47')
// (21, 23, 'sp4_h_r_1')
// (22, 23, 'sp4_h_r_12')
// (23, 23, 'sp4_h_r_25')
// (24, 23, 'sp4_h_r_36')
// (24, 24, 'sp4_r_v_b_43')
// (24, 25, 'sp4_r_v_b_30')
// (24, 26, 'local_g3_3')
// (24, 26, 'lutff_0/in_2')
// (24, 26, 'lutff_1/in_1')
// (24, 26, 'sp4_r_v_b_19')
// (24, 27, 'sp4_r_v_b_6')
// (25, 23, 'sp4_h_l_36')
// (25, 23, 'sp4_v_t_43')
// (25, 24, 'sp4_v_b_43')
// (25, 25, 'sp4_v_b_30')
// (25, 26, 'sp4_v_b_19')
// (25, 27, 'sp4_v_b_6')

wire n59;
// (7, 17, 'sp4_r_v_b_42')
// (7, 18, 'sp4_r_v_b_31')
// (7, 19, 'sp4_r_v_b_18')
// (7, 20, 'sp4_r_v_b_7')
// (7, 21, 'sp4_r_v_b_38')
// (7, 22, 'sp4_r_v_b_27')
// (7, 23, 'sp4_r_v_b_14')
// (7, 24, 'sp4_r_v_b_3')
// (7, 25, 'sp4_r_v_b_43')
// (7, 26, 'sp4_r_v_b_30')
// (7, 27, 'sp4_r_v_b_19')
// (7, 27, 'sp4_r_v_b_43')
// (7, 28, 'sp4_r_v_b_30')
// (7, 28, 'sp4_r_v_b_6')
// (7, 29, 'sp4_r_v_b_19')
// (7, 30, 'sp4_r_v_b_6')
// (8, 16, 'sp4_v_t_42')
// (8, 17, 'sp4_v_b_42')
// (8, 18, 'sp4_v_b_31')
// (8, 19, 'local_g0_2')
// (8, 19, 'ram/RCLKE')
// (8, 19, 'sp4_v_b_18')
// (8, 20, 'sp4_h_r_3')
// (8, 20, 'sp4_h_r_7')
// (8, 20, 'sp4_v_b_7')
// (8, 20, 'sp4_v_t_38')
// (8, 21, 'sp4_v_b_38')
// (8, 22, 'sp4_v_b_27')
// (8, 23, 'sp4_v_b_14')
// (8, 24, 'sp4_v_b_3')
// (8, 24, 'sp4_v_t_43')
// (8, 25, 'sp4_v_b_43')
// (8, 26, 'sp4_v_b_30')
// (8, 26, 'sp4_v_t_43')
// (8, 27, 'local_g1_3')
// (8, 27, 'ram/RCLKE')
// (8, 27, 'sp4_v_b_19')
// (8, 27, 'sp4_v_b_43')
// (8, 28, 'sp4_v_b_30')
// (8, 28, 'sp4_v_b_6')
// (8, 29, 'local_g1_3')
// (8, 29, 'ram/RCLKE')
// (8, 29, 'sp4_v_b_19')
// (8, 30, 'sp4_h_r_6')
// (8, 30, 'sp4_v_b_6')
// (9, 20, 'sp4_h_r_14')
// (9, 20, 'sp4_h_r_18')
// (9, 30, 'sp4_h_r_19')
// (10, 20, 'sp4_h_r_27')
// (10, 20, 'sp4_h_r_31')
// (10, 30, 'sp4_h_r_30')
// (11, 20, 'sp4_h_r_38')
// (11, 20, 'sp4_h_r_42')
// (11, 30, 'sp12_h_r_0')
// (11, 30, 'sp4_h_r_43')
// (12, 20, 'sp4_h_l_38')
// (12, 20, 'sp4_h_l_42')
// (12, 20, 'sp4_h_r_7')
// (12, 30, 'sp12_h_r_3')
// (12, 30, 'sp4_h_l_43')
// (12, 30, 'sp4_h_r_3')
// (13, 20, 'sp4_h_r_18')
// (13, 30, 'sp12_h_r_4')
// (13, 30, 'sp4_h_r_14')
// (14, 20, 'sp4_h_r_31')
// (14, 30, 'sp12_h_r_7')
// (14, 30, 'sp4_h_r_27')
// (15, 20, 'sp4_h_r_42')
// (15, 30, 'sp12_h_r_8')
// (15, 30, 'sp4_h_r_38')
// (16, 20, 'local_g0_4')
// (16, 20, 'lutff_4/in_2')
// (16, 20, 'sp4_h_l_42')
// (16, 20, 'sp4_h_r_4')
// (16, 30, 'sp12_h_r_11')
// (16, 30, 'sp4_h_l_38')
// (17, 20, 'sp4_h_r_17')
// (17, 30, 'sp12_h_r_12')
// (18, 20, 'sp4_h_r_28')
// (18, 30, 'sp12_h_r_15')
// (19, 20, 'sp4_h_r_41')
// (19, 30, 'sp12_h_r_16')
// (20, 20, 'sp4_h_l_41')
// (20, 20, 'sp4_h_r_1')
// (20, 30, 'sp12_h_r_19')
// (21, 20, 'sp4_h_r_12')
// (21, 30, 'sp12_h_r_20')
// (22, 19, 'neigh_op_tnr_2')
// (22, 20, 'neigh_op_rgt_2')
// (22, 20, 'sp4_h_r_25')
// (22, 21, 'neigh_op_bnr_2')
// (22, 30, 'sp12_h_r_23')
// (23, 18, 'sp12_v_t_23')
// (23, 18, 'sp4_r_v_b_45')
// (23, 19, 'neigh_op_top_2')
// (23, 19, 'sp12_v_b_23')
// (23, 19, 'sp4_r_v_b_32')
// (23, 20, 'lutff_2/out')
// (23, 20, 'sp12_v_b_20')
// (23, 20, 'sp4_h_r_36')
// (23, 20, 'sp4_r_v_b_21')
// (23, 21, 'neigh_op_bot_2')
// (23, 21, 'sp12_v_b_19')
// (23, 21, 'sp4_r_v_b_8')
// (23, 22, 'sp12_v_b_16')
// (23, 22, 'sp4_r_v_b_46')
// (23, 23, 'sp12_v_b_15')
// (23, 23, 'sp4_r_v_b_35')
// (23, 24, 'sp12_v_b_12')
// (23, 24, 'sp4_r_v_b_22')
// (23, 25, 'sp12_v_b_11')
// (23, 25, 'sp4_r_v_b_11')
// (23, 26, 'sp12_v_b_8')
// (23, 26, 'sp4_r_v_b_42')
// (23, 27, 'sp12_v_b_7')
// (23, 27, 'sp4_r_v_b_31')
// (23, 28, 'sp12_v_b_4')
// (23, 28, 'sp4_r_v_b_18')
// (23, 29, 'sp12_v_b_3')
// (23, 29, 'sp4_r_v_b_7')
// (23, 30, 'sp12_h_l_23')
// (23, 30, 'sp12_v_b_0')
// (24, 17, 'sp4_v_t_45')
// (24, 18, 'sp4_v_b_45')
// (24, 19, 'neigh_op_tnl_2')
// (24, 19, 'sp4_v_b_32')
// (24, 20, 'neigh_op_lft_2')
// (24, 20, 'sp4_h_l_36')
// (24, 20, 'sp4_v_b_21')
// (24, 21, 'neigh_op_bnl_2')
// (24, 21, 'sp4_v_b_8')
// (24, 21, 'sp4_v_t_46')
// (24, 22, 'sp4_v_b_46')
// (24, 23, 'sp4_v_b_35')
// (24, 24, 'sp4_v_b_22')
// (24, 25, 'sp4_v_b_11')
// (24, 25, 'sp4_v_t_42')
// (24, 26, 'sp4_v_b_42')
// (24, 27, 'sp4_v_b_31')
// (24, 28, 'sp4_v_b_18')
// (24, 29, 'sp4_h_r_7')
// (24, 29, 'sp4_v_b_7')
// (25, 29, 'local_g0_2')
// (25, 29, 'ram/RCLKE')
// (25, 29, 'sp4_h_r_18')
// (26, 29, 'sp4_h_r_31')
// (27, 29, 'sp4_h_r_42')
// (28, 29, 'sp4_h_l_42')

wire n60;
// (7, 18, 'neigh_op_tnr_4')
// (7, 19, 'local_g2_4')
// (7, 19, 'lutff_2/in_2')
// (7, 19, 'neigh_op_rgt_4')
// (7, 20, 'neigh_op_bnr_4')
// (8, 18, 'neigh_op_top_4')
// (8, 19, 'ram/RDATA_11')
// (8, 20, 'neigh_op_bot_4')
// (9, 18, 'neigh_op_tnl_4')
// (9, 19, 'neigh_op_lft_4')
// (9, 20, 'neigh_op_bnl_4')

wire n61;
// (7, 18, 'sp4_r_v_b_46')
// (7, 19, 'sp4_r_v_b_35')
// (7, 20, 'sp4_r_v_b_22')
// (7, 21, 'local_g2_3')
// (7, 21, 'lutff_7/in_2')
// (7, 21, 'sp4_r_v_b_11')
// (8, 17, 'sp4_v_t_46')
// (8, 18, 'sp4_v_b_46')
// (8, 19, 'sp4_v_b_35')
// (8, 20, 'sp4_v_b_22')
// (8, 21, 'sp4_h_r_6')
// (8, 21, 'sp4_v_b_11')
// (9, 21, 'sp4_h_r_19')
// (10, 21, 'sp4_h_r_30')
// (11, 21, 'sp4_h_r_43')
// (12, 21, 'sp4_h_l_43')
// (12, 21, 'sp4_h_r_6')
// (13, 21, 'sp4_h_r_19')
// (14, 21, 'sp4_h_r_30')
// (15, 21, 'sp4_h_r_43')
// (16, 21, 'sp4_h_l_43')
// (16, 21, 'sp4_h_r_6')
// (17, 21, 'sp4_h_r_19')
// (18, 21, 'sp4_h_r_30')
// (19, 21, 'sp4_h_r_43')
// (20, 21, 'sp4_h_l_43')
// (20, 21, 'sp4_h_r_10')
// (21, 21, 'sp4_h_r_23')
// (22, 21, 'sp4_h_r_34')
// (23, 21, 'sp4_h_r_47')
// (23, 22, 'sp4_r_v_b_47')
// (23, 23, 'sp4_r_v_b_34')
// (23, 24, 'neigh_op_tnr_5')
// (23, 24, 'sp4_r_v_b_23')
// (23, 25, 'neigh_op_rgt_5')
// (23, 25, 'sp4_r_v_b_10')
// (23, 26, 'neigh_op_bnr_5')
// (24, 21, 'sp4_h_l_47')
// (24, 21, 'sp4_v_t_47')
// (24, 22, 'sp4_v_b_47')
// (24, 23, 'sp4_v_b_34')
// (24, 24, 'neigh_op_top_5')
// (24, 24, 'sp4_v_b_23')
// (24, 25, 'lutff_5/out')
// (24, 25, 'sp4_v_b_10')
// (24, 26, 'neigh_op_bot_5')
// (25, 24, 'neigh_op_tnl_5')
// (25, 25, 'neigh_op_lft_5')
// (25, 26, 'neigh_op_bnl_5')

wire n62;
// (7, 19, 'local_g1_0')
// (7, 19, 'lutff_3/in_0')
// (7, 19, 'sp4_h_r_8')
// (8, 18, 'neigh_op_tnr_0')
// (8, 19, 'neigh_op_rgt_0')
// (8, 19, 'sp4_h_r_21')
// (8, 20, 'neigh_op_bnr_0')
// (9, 18, 'neigh_op_top_0')
// (9, 19, 'lutff_0/out')
// (9, 19, 'sp4_h_r_32')
// (9, 20, 'neigh_op_bot_0')
// (10, 18, 'neigh_op_tnl_0')
// (10, 19, 'neigh_op_lft_0')
// (10, 19, 'sp4_h_r_45')
// (10, 20, 'neigh_op_bnl_0')
// (11, 19, 'sp4_h_l_45')

wire n63;
// (7, 19, 'local_g1_2')
// (7, 19, 'lutff_0/in_3')
// (7, 19, 'sp4_h_r_10')
// (8, 18, 'neigh_op_tnr_1')
// (8, 19, 'neigh_op_rgt_1')
// (8, 19, 'sp4_h_r_23')
// (8, 20, 'neigh_op_bnr_1')
// (9, 18, 'neigh_op_top_1')
// (9, 19, 'lutff_1/out')
// (9, 19, 'sp4_h_r_34')
// (9, 20, 'neigh_op_bot_1')
// (10, 18, 'neigh_op_tnl_1')
// (10, 19, 'neigh_op_lft_1')
// (10, 19, 'sp4_h_r_47')
// (10, 20, 'neigh_op_bnl_1')
// (11, 19, 'sp4_h_l_47')

wire n64;
// (7, 19, 'neigh_op_tnr_4')
// (7, 20, 'neigh_op_rgt_4')
// (7, 21, 'neigh_op_bnr_4')
// (8, 19, 'neigh_op_top_4')
// (8, 20, 'ram/RDATA_3')
// (8, 21, 'neigh_op_bot_4')
// (9, 19, 'local_g2_4')
// (9, 19, 'lutff_2/in_0')
// (9, 19, 'neigh_op_tnl_4')
// (9, 20, 'neigh_op_lft_4')
// (9, 21, 'neigh_op_bnl_4')

wire n65;
// (7, 19, 'sp4_r_v_b_40')
// (7, 20, 'sp4_r_v_b_29')
// (7, 21, 'local_g3_0')
// (7, 21, 'lutff_5/in_0')
// (7, 21, 'sp4_r_v_b_16')
// (7, 22, 'sp4_r_v_b_5')
// (8, 18, 'sp4_v_t_40')
// (8, 19, 'sp4_v_b_40')
// (8, 20, 'sp4_v_b_29')
// (8, 21, 'sp4_v_b_16')
// (8, 22, 'sp4_h_r_5')
// (8, 22, 'sp4_v_b_5')
// (9, 22, 'sp4_h_r_16')
// (10, 22, 'sp4_h_r_29')
// (11, 22, 'sp4_h_r_40')
// (12, 22, 'sp4_h_l_40')
// (12, 22, 'sp4_h_r_2')
// (13, 22, 'sp4_h_r_15')
// (14, 22, 'sp4_h_r_26')
// (15, 22, 'sp4_h_r_39')
// (16, 22, 'sp4_h_l_39')
// (16, 22, 'sp4_h_r_11')
// (17, 22, 'sp4_h_r_22')
// (18, 22, 'sp4_h_r_35')
// (19, 22, 'sp4_h_r_46')
// (20, 22, 'sp4_h_l_46')
// (20, 22, 'sp4_h_r_3')
// (21, 22, 'sp4_h_r_14')
// (22, 22, 'sp4_h_r_27')
// (23, 22, 'sp4_h_r_38')
// (23, 23, 'sp4_r_v_b_38')
// (23, 24, 'neigh_op_tnr_7')
// (23, 24, 'sp4_r_v_b_27')
// (23, 25, 'neigh_op_rgt_7')
// (23, 25, 'sp4_r_v_b_14')
// (23, 26, 'neigh_op_bnr_7')
// (23, 26, 'sp4_r_v_b_3')
// (24, 22, 'sp4_h_l_38')
// (24, 22, 'sp4_v_t_38')
// (24, 23, 'sp4_v_b_38')
// (24, 24, 'neigh_op_top_7')
// (24, 24, 'sp4_v_b_27')
// (24, 25, 'lutff_7/out')
// (24, 25, 'sp4_v_b_14')
// (24, 26, 'neigh_op_bot_7')
// (24, 26, 'sp4_v_b_3')
// (25, 24, 'neigh_op_tnl_7')
// (25, 25, 'neigh_op_lft_7')
// (25, 26, 'neigh_op_bnl_7')

wire n66;
// (7, 19, 'sp4_r_v_b_43')
// (7, 20, 'sp4_r_v_b_30')
// (7, 21, 'sp4_r_v_b_19')
// (7, 22, 'sp4_r_v_b_6')
// (7, 23, 'sp4_h_r_6')
// (7, 23, 'sp4_r_v_b_43')
// (7, 24, 'sp4_r_v_b_30')
// (7, 25, 'sp4_r_v_b_19')
// (7, 26, 'sp4_r_v_b_6')
// (8, 17, 'local_g3_3')
// (8, 17, 'ram/RCLKE')
// (8, 17, 'sp4_r_v_b_43')
// (8, 18, 'sp4_r_v_b_30')
// (8, 18, 'sp4_v_t_43')
// (8, 19, 'sp4_r_v_b_19')
// (8, 19, 'sp4_v_b_43')
// (8, 20, 'sp4_r_v_b_6')
// (8, 20, 'sp4_v_b_30')
// (8, 21, 'local_g1_3')
// (8, 21, 'ram/RCLKE')
// (8, 21, 'sp4_v_b_19')
// (8, 22, 'sp4_h_r_6')
// (8, 22, 'sp4_v_b_6')
// (8, 22, 'sp4_v_t_43')
// (8, 23, 'local_g1_3')
// (8, 23, 'ram/RCLKE')
// (8, 23, 'sp4_h_r_19')
// (8, 23, 'sp4_v_b_43')
// (8, 24, 'sp4_v_b_30')
// (8, 25, 'local_g1_3')
// (8, 25, 'ram/RCLKE')
// (8, 25, 'sp4_v_b_19')
// (8, 26, 'sp4_v_b_6')
// (9, 16, 'sp4_v_t_43')
// (9, 17, 'sp4_v_b_43')
// (9, 18, 'sp4_v_b_30')
// (9, 19, 'sp4_v_b_19')
// (9, 20, 'sp4_h_r_6')
// (9, 20, 'sp4_v_b_6')
// (9, 22, 'sp4_h_r_19')
// (9, 23, 'sp4_h_r_30')
// (10, 20, 'sp4_h_r_19')
// (10, 22, 'sp4_h_r_30')
// (10, 23, 'sp4_h_r_43')
// (11, 20, 'sp4_h_r_30')
// (11, 22, 'sp4_h_r_43')
// (11, 23, 'sp4_h_l_43')
// (11, 23, 'sp4_h_r_10')
// (12, 20, 'sp4_h_r_43')
// (12, 22, 'sp4_h_l_43')
// (12, 22, 'sp4_h_r_6')
// (12, 23, 'sp4_h_r_23')
// (13, 20, 'sp4_h_l_43')
// (13, 20, 'sp4_h_r_6')
// (13, 22, 'sp4_h_r_19')
// (13, 23, 'sp4_h_r_34')
// (14, 20, 'sp4_h_r_19')
// (14, 22, 'sp4_h_r_30')
// (14, 23, 'sp4_h_r_47')
// (15, 20, 'sp4_h_r_30')
// (15, 22, 'sp4_h_r_43')
// (15, 23, 'sp4_h_l_47')
// (15, 23, 'sp4_h_r_10')
// (16, 20, 'sp4_h_r_43')
// (16, 22, 'sp4_h_l_43')
// (16, 22, 'sp4_h_r_6')
// (16, 23, 'sp4_h_r_23')
// (17, 20, 'sp4_h_l_43')
// (17, 20, 'sp4_h_r_3')
// (17, 22, 'sp4_h_r_19')
// (17, 23, 'sp4_h_r_34')
// (18, 20, 'sp4_h_r_14')
// (18, 22, 'sp4_h_r_30')
// (18, 23, 'sp4_h_r_47')
// (19, 20, 'sp4_h_r_27')
// (19, 22, 'sp4_h_r_43')
// (19, 23, 'sp4_h_l_47')
// (19, 23, 'sp4_h_r_10')
// (20, 20, 'sp4_h_r_38')
// (20, 22, 'sp4_h_l_43')
// (20, 22, 'sp4_h_r_6')
// (20, 23, 'sp4_h_r_23')
// (21, 20, 'sp4_h_l_38')
// (21, 20, 'sp4_h_r_0')
// (21, 22, 'sp4_h_r_19')
// (21, 23, 'sp4_h_r_34')
// (22, 19, 'neigh_op_tnr_4')
// (22, 20, 'neigh_op_rgt_4')
// (22, 20, 'sp4_h_r_13')
// (22, 20, 'sp4_r_v_b_40')
// (22, 21, 'neigh_op_bnr_4')
// (22, 21, 'sp4_r_v_b_29')
// (22, 22, 'sp4_h_r_30')
// (22, 22, 'sp4_r_v_b_16')
// (22, 23, 'sp4_h_r_47')
// (22, 23, 'sp4_r_v_b_5')
// (23, 19, 'neigh_op_top_4')
// (23, 19, 'sp4_r_v_b_36')
// (23, 19, 'sp4_v_t_40')
// (23, 20, 'lutff_4/out')
// (23, 20, 'sp4_h_r_24')
// (23, 20, 'sp4_r_v_b_25')
// (23, 20, 'sp4_v_b_40')
// (23, 21, 'neigh_op_bot_4')
// (23, 21, 'sp4_r_v_b_12')
// (23, 21, 'sp4_v_b_29')
// (23, 22, 'sp4_h_r_43')
// (23, 22, 'sp4_r_v_b_1')
// (23, 22, 'sp4_v_b_16')
// (23, 23, 'sp4_h_l_47')
// (23, 23, 'sp4_v_b_5')
// (24, 18, 'sp4_v_t_36')
// (24, 19, 'neigh_op_tnl_4')
// (24, 19, 'sp4_v_b_36')
// (24, 20, 'neigh_op_lft_4')
// (24, 20, 'sp4_h_r_37')
// (24, 20, 'sp4_v_b_25')
// (24, 21, 'neigh_op_bnl_4')
// (24, 21, 'sp4_v_b_12')
// (24, 22, 'sp4_h_l_43')
// (24, 22, 'sp4_v_b_1')
// (25, 20, 'sp4_h_l_37')

wire n67;
// (7, 20, 'lutff_1/cout')
// (7, 20, 'lutff_2/in_3')

wire n68;
// (7, 20, 'lutff_2/cout')
// (7, 20, 'lutff_3/in_3')

wire n69;
// (7, 20, 'lutff_3/cout')
// (7, 20, 'lutff_4/in_3')

wire n70;
// (7, 20, 'lutff_4/cout')
// (7, 20, 'lutff_5/in_3')

wire n71;
// (7, 20, 'lutff_5/cout')
// (7, 20, 'lutff_6/in_3')

wire n72;
// (7, 20, 'lutff_6/cout')
// (7, 20, 'lutff_7/in_3')

wire n73;
// (7, 20, 'neigh_op_tnr_4')
// (7, 21, 'local_g2_4')
// (7, 21, 'lutff_6/in_0')
// (7, 21, 'neigh_op_rgt_4')
// (7, 22, 'neigh_op_bnr_4')
// (8, 20, 'neigh_op_top_4')
// (8, 21, 'ram/RDATA_11')
// (8, 22, 'neigh_op_bot_4')
// (9, 20, 'neigh_op_tnl_4')
// (9, 21, 'neigh_op_lft_4')
// (9, 22, 'neigh_op_bnl_4')

wire n74;
// (7, 21, 'local_g3_4')
// (7, 21, 'lutff_2/in_3')
// (7, 21, 'neigh_op_tnr_4')
// (7, 22, 'neigh_op_rgt_4')
// (7, 23, 'neigh_op_bnr_4')
// (8, 21, 'neigh_op_top_4')
// (8, 22, 'ram/RDATA_3')
// (8, 23, 'neigh_op_bot_4')
// (9, 21, 'neigh_op_tnl_4')
// (9, 22, 'neigh_op_lft_4')
// (9, 23, 'neigh_op_bnl_4')

wire n75;
// (7, 21, 'sp4_r_v_b_42')
// (7, 22, 'sp4_r_v_b_31')
// (7, 23, 'local_g3_2')
// (7, 23, 'lutff_5/in_2')
// (7, 23, 'sp4_r_v_b_18')
// (7, 24, 'sp4_r_v_b_7')
// (8, 20, 'sp4_h_r_1')
// (8, 20, 'sp4_v_t_42')
// (8, 21, 'sp4_v_b_42')
// (8, 22, 'sp4_v_b_31')
// (8, 23, 'sp4_v_b_18')
// (8, 24, 'sp4_v_b_7')
// (9, 20, 'sp4_h_r_12')
// (10, 20, 'sp4_h_r_25')
// (11, 20, 'sp4_h_r_36')
// (12, 20, 'sp4_h_l_36')
// (12, 20, 'sp4_h_r_10')
// (13, 20, 'sp4_h_r_23')
// (14, 20, 'sp4_h_r_34')
// (15, 20, 'sp4_h_r_47')
// (16, 20, 'sp4_h_l_47')
// (16, 20, 'sp4_h_r_7')
// (17, 20, 'sp4_h_r_18')
// (18, 20, 'sp4_h_r_31')
// (19, 20, 'sp4_h_r_42')
// (20, 20, 'sp4_h_l_42')
// (20, 20, 'sp4_h_r_11')
// (21, 20, 'sp4_h_r_22')
// (22, 20, 'sp4_h_r_35')
// (23, 16, 'neigh_op_tnr_7')
// (23, 17, 'neigh_op_rgt_7')
// (23, 17, 'sp4_r_v_b_46')
// (23, 18, 'neigh_op_bnr_7')
// (23, 18, 'sp4_r_v_b_35')
// (23, 19, 'sp4_r_v_b_22')
// (23, 20, 'sp4_h_r_46')
// (23, 20, 'sp4_r_v_b_11')
// (24, 16, 'neigh_op_top_7')
// (24, 16, 'sp4_v_t_46')
// (24, 17, 'lutff_7/out')
// (24, 17, 'sp4_v_b_46')
// (24, 18, 'neigh_op_bot_7')
// (24, 18, 'sp4_v_b_35')
// (24, 19, 'sp4_v_b_22')
// (24, 20, 'sp4_h_l_46')
// (24, 20, 'sp4_v_b_11')
// (25, 16, 'neigh_op_tnl_7')
// (25, 17, 'neigh_op_lft_7')
// (25, 18, 'neigh_op_bnl_7')

wire n76;
// (7, 22, 'neigh_op_tnr_4')
// (7, 23, 'local_g2_4')
// (7, 23, 'lutff_0/in_0')
// (7, 23, 'neigh_op_rgt_4')
// (7, 24, 'neigh_op_bnr_4')
// (8, 22, 'neigh_op_top_4')
// (8, 23, 'ram/RDATA_11')
// (8, 24, 'neigh_op_bot_4')
// (9, 22, 'neigh_op_tnl_4')
// (9, 23, 'neigh_op_lft_4')
// (9, 24, 'neigh_op_bnl_4')

wire n77;
// (7, 22, 'sp4_r_v_b_45')
// (7, 23, 'local_g0_3')
// (7, 23, 'lutff_0/in_1')
// (7, 23, 'sp4_r_v_b_32')
// (7, 24, 'sp4_r_v_b_21')
// (7, 25, 'sp4_r_v_b_8')
// (7, 26, 'sp4_r_v_b_45')
// (7, 27, 'sp4_r_v_b_32')
// (7, 28, 'neigh_op_tnr_4')
// (7, 28, 'sp4_r_v_b_21')
// (7, 29, 'neigh_op_rgt_4')
// (7, 29, 'sp4_r_v_b_8')
// (7, 30, 'neigh_op_bnr_4')
// (8, 21, 'sp4_v_t_45')
// (8, 22, 'sp4_v_b_45')
// (8, 23, 'sp4_v_b_32')
// (8, 24, 'sp4_v_b_21')
// (8, 25, 'sp4_v_b_8')
// (8, 25, 'sp4_v_t_45')
// (8, 26, 'sp4_v_b_45')
// (8, 27, 'sp4_v_b_32')
// (8, 28, 'neigh_op_top_4')
// (8, 28, 'sp4_v_b_21')
// (8, 29, 'ram/RDATA_11')
// (8, 29, 'sp4_v_b_8')
// (8, 30, 'neigh_op_bot_4')
// (9, 28, 'neigh_op_tnl_4')
// (9, 29, 'neigh_op_lft_4')
// (9, 30, 'neigh_op_bnl_4')

wire n78;
// (7, 23, 'local_g3_4')
// (7, 23, 'lutff_6/in_1')
// (7, 23, 'neigh_op_tnr_4')
// (7, 24, 'neigh_op_rgt_4')
// (7, 25, 'neigh_op_bnr_4')
// (8, 23, 'neigh_op_top_4')
// (8, 24, 'ram/RDATA_3')
// (8, 25, 'neigh_op_bot_4')
// (9, 23, 'neigh_op_tnl_4')
// (9, 24, 'neigh_op_lft_4')
// (9, 25, 'neigh_op_bnl_4')

wire n79;
// (7, 23, 'local_g3_5')
// (7, 23, 'lutff_5/in_1')
// (7, 23, 'sp4_r_v_b_45')
// (7, 24, 'sp4_r_v_b_32')
// (7, 25, 'sp4_r_v_b_21')
// (7, 26, 'sp4_r_v_b_8')
// (7, 27, 'sp4_r_v_b_45')
// (7, 28, 'sp4_r_v_b_32')
// (7, 29, 'neigh_op_tnr_4')
// (7, 29, 'sp4_r_v_b_21')
// (7, 30, 'neigh_op_rgt_4')
// (7, 30, 'sp4_r_v_b_8')
// (7, 31, 'neigh_op_bnr_4')
// (8, 22, 'sp4_v_t_45')
// (8, 23, 'sp4_v_b_45')
// (8, 24, 'sp4_v_b_32')
// (8, 25, 'sp4_v_b_21')
// (8, 26, 'sp4_v_b_8')
// (8, 26, 'sp4_v_t_45')
// (8, 27, 'sp4_v_b_45')
// (8, 28, 'sp4_v_b_32')
// (8, 29, 'neigh_op_top_4')
// (8, 29, 'sp4_v_b_21')
// (8, 30, 'ram/RDATA_3')
// (8, 30, 'sp4_v_b_8')
// (8, 31, 'neigh_op_bot_4')
// (9, 29, 'neigh_op_tnl_4')
// (9, 30, 'neigh_op_lft_4')
// (9, 31, 'neigh_op_bnl_4')

reg n80 = 0;
// (7, 23, 'sp12_h_r_1')
// (8, 23, 'sp12_h_r_2')
// (9, 17, 'sp4_r_v_b_46')
// (9, 18, 'sp4_r_v_b_35')
// (9, 19, 'local_g3_6')
// (9, 19, 'lutff_0/in_3')
// (9, 19, 'lutff_1/in_0')
// (9, 19, 'sp4_r_v_b_22')
// (9, 20, 'sp4_r_v_b_11')
// (9, 23, 'local_g1_5')
// (9, 23, 'lutff_3/in_3')
// (9, 23, 'sp12_h_r_5')
// (10, 16, 'sp4_v_t_46')
// (10, 17, 'sp4_v_b_46')
// (10, 18, 'sp4_v_b_35')
// (10, 19, 'sp4_v_b_22')
// (10, 20, 'sp4_h_r_6')
// (10, 20, 'sp4_v_b_11')
// (10, 23, 'sp12_h_r_6')
// (11, 20, 'sp4_h_r_19')
// (11, 23, 'sp12_h_r_9')
// (12, 20, 'sp4_h_r_30')
// (12, 23, 'sp12_h_r_10')
// (13, 20, 'sp4_h_r_43')
// (13, 23, 'sp12_h_r_13')
// (14, 20, 'sp4_h_l_43')
// (14, 20, 'sp4_h_r_3')
// (14, 23, 'sp12_h_r_14')
// (15, 20, 'sp4_h_r_14')
// (15, 23, 'sp12_h_r_17')
// (16, 20, 'sp4_h_r_27')
// (16, 23, 'sp12_h_r_18')
// (17, 20, 'sp4_h_r_38')
// (17, 21, 'sp4_r_v_b_38')
// (17, 22, 'neigh_op_tnr_7')
// (17, 22, 'sp4_r_v_b_27')
// (17, 23, 'neigh_op_rgt_7')
// (17, 23, 'sp12_h_r_21')
// (17, 23, 'sp4_h_r_3')
// (17, 23, 'sp4_r_v_b_14')
// (17, 24, 'neigh_op_bnr_7')
// (17, 24, 'sp4_r_v_b_3')
// (18, 20, 'sp4_h_l_38')
// (18, 20, 'sp4_v_t_38')
// (18, 21, 'sp4_v_b_38')
// (18, 22, 'neigh_op_top_7')
// (18, 22, 'sp4_r_v_b_42')
// (18, 22, 'sp4_v_b_27')
// (18, 23, 'lutff_7/out')
// (18, 23, 'sp12_h_r_22')
// (18, 23, 'sp4_h_r_14')
// (18, 23, 'sp4_r_v_b_31')
// (18, 23, 'sp4_v_b_14')
// (18, 24, 'neigh_op_bot_7')
// (18, 24, 'sp4_r_v_b_18')
// (18, 24, 'sp4_v_b_3')
// (18, 25, 'sp4_r_v_b_7')
// (19, 21, 'sp4_h_r_0')
// (19, 21, 'sp4_v_t_42')
// (19, 22, 'neigh_op_tnl_7')
// (19, 22, 'sp4_v_b_42')
// (19, 23, 'neigh_op_lft_7')
// (19, 23, 'sp12_h_l_22')
// (19, 23, 'sp4_h_r_27')
// (19, 23, 'sp4_v_b_31')
// (19, 24, 'neigh_op_bnl_7')
// (19, 24, 'sp4_v_b_18')
// (19, 25, 'sp4_h_r_1')
// (19, 25, 'sp4_v_b_7')
// (20, 21, 'sp4_h_r_13')
// (20, 23, 'sp4_h_r_38')
// (20, 25, 'sp4_h_r_12')
// (21, 21, 'sp4_h_r_24')
// (21, 23, 'sp4_h_l_38')
// (21, 23, 'sp4_h_r_3')
// (21, 25, 'sp4_h_r_25')
// (22, 18, 'sp4_r_v_b_37')
// (22, 19, 'sp4_r_v_b_24')
// (22, 20, 'sp4_r_v_b_13')
// (22, 21, 'sp4_h_r_37')
// (22, 21, 'sp4_r_v_b_0')
// (22, 23, 'sp4_h_r_14')
// (22, 25, 'sp4_h_r_36')
// (23, 17, 'sp4_h_r_0')
// (23, 17, 'sp4_v_t_37')
// (23, 18, 'sp4_v_b_37')
// (23, 19, 'sp4_v_b_24')
// (23, 20, 'sp4_v_b_13')
// (23, 21, 'sp4_h_l_37')
// (23, 21, 'sp4_h_r_3')
// (23, 21, 'sp4_v_b_0')
// (23, 23, 'sp4_h_r_27')
// (23, 25, 'sp4_h_l_36')
// (23, 25, 'sp4_h_r_1')
// (24, 17, 'local_g0_5')
// (24, 17, 'lutff_5/in_0')
// (24, 17, 'lutff_7/in_2')
// (24, 17, 'sp4_h_r_13')
// (24, 20, 'sp4_r_v_b_38')
// (24, 21, 'local_g0_6')
// (24, 21, 'lutff_7/in_1')
// (24, 21, 'sp4_h_r_14')
// (24, 21, 'sp4_r_v_b_27')
// (24, 22, 'local_g2_6')
// (24, 22, 'lutff_7/in_3')
// (24, 22, 'sp4_r_v_b_14')
// (24, 23, 'sp4_h_r_38')
// (24, 23, 'sp4_r_v_b_3')
// (24, 25, 'local_g0_4')
// (24, 25, 'lutff_5/in_1')
// (24, 25, 'lutff_7/in_1')
// (24, 25, 'sp4_h_r_12')
// (25, 17, 'sp4_h_r_24')
// (25, 19, 'sp4_v_t_38')
// (25, 20, 'sp4_v_b_38')
// (25, 21, 'sp4_h_r_27')
// (25, 21, 'sp4_v_b_27')
// (25, 22, 'sp4_v_b_14')
// (25, 23, 'sp4_h_l_38')
// (25, 23, 'sp4_v_b_3')
// (25, 25, 'sp4_h_r_25')
// (26, 17, 'sp4_h_r_37')
// (26, 21, 'sp4_h_r_38')
// (26, 25, 'sp4_h_r_36')
// (27, 17, 'sp4_h_l_37')
// (27, 21, 'sp4_h_l_38')
// (27, 25, 'sp4_h_l_36')

wire n81;
// (7, 24, 'neigh_op_tnr_4')
// (7, 25, 'local_g3_4')
// (7, 25, 'lutff_0/in_3')
// (7, 25, 'neigh_op_rgt_4')
// (7, 26, 'neigh_op_bnr_4')
// (8, 24, 'neigh_op_top_4')
// (8, 25, 'ram/RDATA_11')
// (8, 26, 'neigh_op_bot_4')
// (9, 24, 'neigh_op_tnl_4')
// (9, 25, 'neigh_op_lft_4')
// (9, 26, 'neigh_op_bnl_4')

wire n82;
// (7, 24, 'sp4_r_v_b_45')
// (7, 25, 'local_g2_0')
// (7, 25, 'lutff_0/in_0')
// (7, 25, 'sp4_r_v_b_32')
// (7, 26, 'neigh_op_tnr_4')
// (7, 26, 'sp4_r_v_b_21')
// (7, 27, 'neigh_op_rgt_4')
// (7, 27, 'sp4_r_v_b_8')
// (7, 28, 'neigh_op_bnr_4')
// (8, 23, 'sp4_v_t_45')
// (8, 24, 'sp4_v_b_45')
// (8, 25, 'sp4_v_b_32')
// (8, 26, 'neigh_op_top_4')
// (8, 26, 'sp4_v_b_21')
// (8, 27, 'ram/RDATA_11')
// (8, 27, 'sp4_v_b_8')
// (8, 28, 'neigh_op_bot_4')
// (9, 26, 'neigh_op_tnl_4')
// (9, 27, 'neigh_op_lft_4')
// (9, 28, 'neigh_op_bnl_4')

wire n83;
// (7, 25, 'neigh_op_tnr_4')
// (7, 26, 'neigh_op_rgt_4')
// (7, 27, 'neigh_op_bnr_4')
// (8, 25, 'neigh_op_top_4')
// (8, 26, 'ram/RDATA_3')
// (8, 27, 'neigh_op_bot_4')
// (9, 25, 'local_g2_4')
// (9, 25, 'lutff_6/in_2')
// (9, 25, 'neigh_op_tnl_4')
// (9, 26, 'neigh_op_lft_4')
// (9, 27, 'neigh_op_bnl_4')

wire n84;
// (7, 27, 'neigh_op_tnr_4')
// (7, 28, 'neigh_op_rgt_4')
// (7, 29, 'neigh_op_bnr_4')
// (8, 25, 'sp4_r_v_b_44')
// (8, 26, 'sp4_r_v_b_33')
// (8, 27, 'neigh_op_top_4')
// (8, 27, 'sp4_r_v_b_20')
// (8, 28, 'ram/RDATA_3')
// (8, 28, 'sp4_r_v_b_9')
// (8, 29, 'neigh_op_bot_4')
// (9, 24, 'sp4_v_t_44')
// (9, 25, 'local_g3_4')
// (9, 25, 'lutff_6/in_3')
// (9, 25, 'sp4_v_b_44')
// (9, 26, 'sp4_v_b_33')
// (9, 27, 'neigh_op_tnl_4')
// (9, 27, 'sp4_v_b_20')
// (9, 28, 'neigh_op_lft_4')
// (9, 28, 'sp4_v_b_9')
// (9, 29, 'neigh_op_bnl_4')

wire n85;
// (8, 18, 'neigh_op_tnr_2')
// (8, 19, 'neigh_op_rgt_2')
// (8, 20, 'neigh_op_bnr_2')
// (9, 18, 'neigh_op_top_2')
// (9, 19, 'local_g0_2')
// (9, 19, 'lutff_1/in_1')
// (9, 19, 'lutff_2/out')
// (9, 20, 'neigh_op_bot_2')
// (10, 18, 'neigh_op_tnl_2')
// (10, 19, 'neigh_op_lft_2')
// (10, 20, 'neigh_op_bnl_2')

reg n86 = 0;
// (8, 19, 'sp4_r_v_b_41')
// (8, 20, 'sp4_r_v_b_28')
// (8, 21, 'sp4_r_v_b_17')
// (8, 22, 'sp4_r_v_b_4')
// (8, 23, 'sp4_r_v_b_41')
// (8, 24, 'sp4_r_v_b_28')
// (8, 25, 'sp4_r_v_b_17')
// (8, 26, 'sp4_r_v_b_4')
// (9, 18, 'sp4_v_t_41')
// (9, 19, 'local_g3_1')
// (9, 19, 'lutff_0/in_2')
// (9, 19, 'lutff_2/in_2')
// (9, 19, 'sp4_v_b_41')
// (9, 20, 'sp4_v_b_28')
// (9, 21, 'sp4_v_b_17')
// (9, 22, 'sp4_h_r_4')
// (9, 22, 'sp4_v_b_4')
// (9, 22, 'sp4_v_t_41')
// (9, 23, 'local_g2_1')
// (9, 23, 'lutff_3/in_2')
// (9, 23, 'sp4_v_b_41')
// (9, 24, 'sp4_v_b_28')
// (9, 25, 'sp4_v_b_17')
// (9, 26, 'sp4_v_b_4')
// (10, 22, 'sp4_h_r_17')
// (11, 22, 'sp4_h_r_28')
// (12, 22, 'sp4_h_r_41')
// (13, 22, 'sp4_h_l_41')
// (13, 22, 'sp4_h_r_1')
// (14, 22, 'sp4_h_r_12')
// (15, 22, 'sp4_h_r_25')
// (16, 22, 'sp4_h_r_36')
// (17, 22, 'sp4_h_l_36')
// (17, 22, 'sp4_h_r_10')
// (18, 22, 'sp4_h_r_23')
// (19, 22, 'sp4_h_r_34')
// (20, 22, 'sp4_h_r_47')
// (21, 22, 'sp4_h_l_47')
// (21, 22, 'sp4_h_r_7')
// (22, 22, 'sp4_h_r_18')
// (23, 15, 'sp4_r_v_b_43')
// (23, 16, 'sp4_r_v_b_30')
// (23, 17, 'sp4_r_v_b_19')
// (23, 18, 'sp4_r_v_b_6')
// (23, 19, 'sp4_r_v_b_47')
// (23, 20, 'sp4_r_v_b_34')
// (23, 21, 'neigh_op_tnr_5')
// (23, 21, 'sp4_r_v_b_23')
// (23, 22, 'neigh_op_rgt_5')
// (23, 22, 'sp4_h_r_31')
// (23, 22, 'sp4_r_v_b_10')
// (23, 23, 'neigh_op_bnr_5')
// (24, 14, 'sp4_v_t_43')
// (24, 15, 'sp12_v_t_22')
// (24, 15, 'sp4_v_b_43')
// (24, 16, 'sp12_v_b_22')
// (24, 16, 'sp4_v_b_30')
// (24, 17, 'local_g1_3')
// (24, 17, 'lutff_5/in_1')
// (24, 17, 'lutff_7/in_1')
// (24, 17, 'sp12_v_b_21')
// (24, 17, 'sp4_v_b_19')
// (24, 18, 'sp12_v_b_18')
// (24, 18, 'sp4_v_b_6')
// (24, 18, 'sp4_v_t_47')
// (24, 19, 'sp12_v_b_17')
// (24, 19, 'sp4_v_b_47')
// (24, 20, 'sp12_v_b_14')
// (24, 20, 'sp4_v_b_34')
// (24, 21, 'local_g1_5')
// (24, 21, 'lutff_7/in_3')
// (24, 21, 'neigh_op_top_5')
// (24, 21, 'sp12_v_b_13')
// (24, 21, 'sp4_v_b_23')
// (24, 22, 'local_g0_5')
// (24, 22, 'lutff_5/out')
// (24, 22, 'lutff_7/in_0')
// (24, 22, 'sp12_v_b_10')
// (24, 22, 'sp4_h_r_42')
// (24, 22, 'sp4_v_b_10')
// (24, 23, 'neigh_op_bot_5')
// (24, 23, 'sp12_v_b_9')
// (24, 24, 'sp12_v_b_6')
// (24, 25, 'sp12_v_b_5')
// (24, 26, 'local_g3_2')
// (24, 26, 'lutff_0/in_1')
// (24, 26, 'lutff_1/in_2')
// (24, 26, 'sp12_v_b_2')
// (24, 27, 'sp12_v_b_1')
// (25, 21, 'neigh_op_tnl_5')
// (25, 22, 'neigh_op_lft_5')
// (25, 22, 'sp4_h_l_42')
// (25, 23, 'neigh_op_bnl_5')

wire n87;
// (9, 17, 'sp4_r_v_b_40')
// (9, 18, 'sp4_r_v_b_29')
// (9, 19, 'local_g3_0')
// (9, 19, 'lutff_2/in_3')
// (9, 19, 'sp4_r_v_b_16')
// (9, 20, 'sp4_r_v_b_5')
// (10, 16, 'sp4_v_t_40')
// (10, 17, 'sp4_v_b_40')
// (10, 18, 'sp4_v_b_29')
// (10, 19, 'sp4_v_b_16')
// (10, 20, 'sp4_h_r_0')
// (10, 20, 'sp4_v_b_5')
// (11, 20, 'sp4_h_r_13')
// (12, 20, 'sp4_h_r_24')
// (13, 20, 'sp4_h_r_37')
// (14, 20, 'sp4_h_l_37')
// (14, 20, 'sp4_h_r_4')
// (15, 20, 'sp4_h_r_17')
// (16, 20, 'sp4_h_r_28')
// (17, 20, 'sp4_h_r_41')
// (18, 20, 'sp4_h_l_41')
// (18, 20, 'sp4_h_r_1')
// (19, 20, 'sp4_h_r_12')
// (20, 20, 'sp4_h_r_25')
// (21, 20, 'sp4_h_r_36')
// (22, 20, 'sp4_h_l_36')
// (22, 20, 'sp4_h_r_5')
// (23, 20, 'sp4_h_r_16')
// (24, 19, 'neigh_op_tnr_4')
// (24, 20, 'neigh_op_rgt_4')
// (24, 20, 'sp4_h_r_29')
// (24, 21, 'neigh_op_bnr_4')
// (25, 19, 'neigh_op_top_4')
// (25, 20, 'ram/RDATA_3')
// (25, 20, 'sp4_h_r_40')
// (25, 21, 'neigh_op_bot_4')
// (26, 19, 'neigh_op_tnl_4')
// (26, 20, 'neigh_op_lft_4')
// (26, 20, 'sp4_h_l_40')
// (26, 21, 'neigh_op_bnl_4')

wire n88;
// (13, 13, 'sp4_h_r_6')
// (14, 13, 'sp4_h_r_19')
// (15, 13, 'neigh_op_tnr_5')
// (15, 13, 'sp4_h_r_30')
// (15, 14, 'neigh_op_rgt_5')
// (15, 15, 'neigh_op_bnr_5')
// (16, 13, 'local_g3_3')
// (16, 13, 'lutff_global/cen')
// (16, 13, 'neigh_op_top_5')
// (16, 13, 'sp4_h_r_43')
// (16, 14, 'lutff_5/out')
// (16, 14, 'sp4_r_v_b_43')
// (16, 15, 'neigh_op_bot_5')
// (16, 15, 'sp4_r_v_b_30')
// (16, 16, 'sp4_r_v_b_19')
// (16, 17, 'sp4_r_v_b_6')
// (17, 13, 'neigh_op_tnl_5')
// (17, 13, 'sp4_h_l_43')
// (17, 13, 'sp4_v_t_43')
// (17, 14, 'neigh_op_lft_5')
// (17, 14, 'sp4_v_b_43')
// (17, 15, 'neigh_op_bnl_5')
// (17, 15, 'sp4_v_b_30')
// (17, 16, 'sp4_v_b_19')
// (17, 17, 'sp4_v_b_6')

reg n89 = 0;
// (14, 14, 'neigh_op_tnr_4')
// (14, 15, 'neigh_op_rgt_4')
// (14, 16, 'neigh_op_bnr_4')
// (15, 14, 'neigh_op_top_4')
// (15, 15, 'lutff_4/out')
// (15, 16, 'neigh_op_bot_4')
// (16, 14, 'local_g3_4')
// (16, 14, 'lutff_4/in_1')
// (16, 14, 'neigh_op_tnl_4')
// (16, 15, 'neigh_op_lft_4')
// (16, 16, 'neigh_op_bnl_4')

reg n90 = 0;
// (14, 14, 'neigh_op_tnr_5')
// (14, 15, 'neigh_op_rgt_5')
// (14, 16, 'neigh_op_bnr_5')
// (15, 14, 'neigh_op_top_5')
// (15, 15, 'local_g3_5')
// (15, 15, 'lutff_4/in_0')
// (15, 15, 'lutff_5/out')
// (15, 16, 'neigh_op_bot_5')
// (16, 14, 'neigh_op_tnl_5')
// (16, 15, 'neigh_op_lft_5')
// (16, 16, 'neigh_op_bnl_5')

reg n91 = 0;
// (15, 10, 'neigh_op_tnr_2')
// (15, 11, 'neigh_op_rgt_2')
// (15, 12, 'neigh_op_bnr_2')
// (16, 10, 'neigh_op_top_2')
// (16, 11, 'local_g3_2')
// (16, 11, 'lutff_2/in_1')
// (16, 11, 'lutff_2/out')
// (16, 12, 'neigh_op_bot_2')
// (17, 10, 'local_g2_2')
// (17, 10, 'lutff_2/in_0')
// (17, 10, 'neigh_op_tnl_2')
// (17, 11, 'local_g0_2')
// (17, 11, 'lutff_3/in_1')
// (17, 11, 'neigh_op_lft_2')
// (17, 12, 'neigh_op_bnl_2')

reg n92 = 0;
// (15, 10, 'neigh_op_tnr_3')
// (15, 11, 'neigh_op_rgt_3')
// (15, 12, 'neigh_op_bnr_3')
// (16, 10, 'neigh_op_top_3')
// (16, 11, 'local_g1_3')
// (16, 11, 'lutff_3/in_1')
// (16, 11, 'lutff_3/out')
// (16, 12, 'neigh_op_bot_3')
// (17, 10, 'neigh_op_tnl_3')
// (17, 11, 'local_g0_3')
// (17, 11, 'lutff_3/in_0')
// (17, 11, 'lutff_4/in_3')
// (17, 11, 'neigh_op_lft_3')
// (17, 12, 'neigh_op_bnl_3')

reg n93 = 0;
// (15, 10, 'neigh_op_tnr_4')
// (15, 11, 'neigh_op_rgt_4')
// (15, 12, 'neigh_op_bnr_4')
// (16, 10, 'neigh_op_top_4')
// (16, 11, 'local_g3_4')
// (16, 11, 'lutff_4/in_1')
// (16, 11, 'lutff_4/out')
// (16, 12, 'neigh_op_bot_4')
// (17, 10, 'local_g3_4')
// (17, 10, 'lutff_3/in_0')
// (17, 10, 'neigh_op_tnl_4')
// (17, 11, 'local_g0_4')
// (17, 11, 'lutff_2/in_2')
// (17, 11, 'neigh_op_lft_4')
// (17, 12, 'neigh_op_bnl_4')

reg n94 = 0;
// (15, 10, 'neigh_op_tnr_5')
// (15, 11, 'neigh_op_rgt_5')
// (15, 12, 'neigh_op_bnr_5')
// (16, 10, 'neigh_op_top_5')
// (16, 11, 'local_g0_5')
// (16, 11, 'lutff_5/in_2')
// (16, 11, 'lutff_5/out')
// (16, 12, 'neigh_op_bot_5')
// (17, 10, 'neigh_op_tnl_5')
// (17, 11, 'local_g0_5')
// (17, 11, 'lutff_1/in_0')
// (17, 11, 'lutff_2/in_1')
// (17, 11, 'neigh_op_lft_5')
// (17, 12, 'neigh_op_bnl_5')

reg n95 = 0;
// (15, 10, 'neigh_op_tnr_6')
// (15, 11, 'neigh_op_rgt_6')
// (15, 12, 'neigh_op_bnr_6')
// (16, 10, 'neigh_op_top_6')
// (16, 11, 'local_g1_6')
// (16, 11, 'lutff_6/in_1')
// (16, 11, 'lutff_6/out')
// (16, 12, 'neigh_op_bot_6')
// (17, 10, 'neigh_op_tnl_6')
// (17, 11, 'local_g0_6')
// (17, 11, 'local_g1_6')
// (17, 11, 'lutff_0/in_3')
// (17, 11, 'lutff_2/in_0')
// (17, 11, 'neigh_op_lft_6')
// (17, 12, 'neigh_op_bnl_6')

reg n96 = 0;
// (15, 10, 'neigh_op_tnr_7')
// (15, 11, 'neigh_op_rgt_7')
// (15, 12, 'neigh_op_bnr_7')
// (16, 10, 'neigh_op_top_7')
// (16, 11, 'local_g1_7')
// (16, 11, 'lutff_7/in_1')
// (16, 11, 'lutff_7/out')
// (16, 12, 'neigh_op_bot_7')
// (17, 10, 'neigh_op_tnl_7')
// (17, 11, 'local_g0_7')
// (17, 11, 'lutff_2/in_3')
// (17, 11, 'lutff_5/in_2')
// (17, 11, 'neigh_op_lft_7')
// (17, 12, 'neigh_op_bnl_7')

reg n97 = 0;
// (15, 11, 'neigh_op_tnr_0')
// (15, 12, 'neigh_op_rgt_0')
// (15, 13, 'neigh_op_bnr_0')
// (16, 11, 'neigh_op_top_0')
// (16, 12, 'local_g2_0')
// (16, 12, 'lutff_0/in_2')
// (16, 12, 'lutff_0/out')
// (16, 13, 'neigh_op_bot_0')
// (17, 11, 'neigh_op_tnl_0')
// (17, 12, 'local_g0_0')
// (17, 12, 'lutff_6/in_0')
// (17, 12, 'neigh_op_lft_0')
// (17, 13, 'local_g3_0')
// (17, 13, 'lutff_7/in_2')
// (17, 13, 'neigh_op_bnl_0')

reg n98 = 0;
// (15, 11, 'neigh_op_tnr_1')
// (15, 12, 'neigh_op_rgt_1')
// (15, 13, 'neigh_op_bnr_1')
// (16, 11, 'neigh_op_top_1')
// (16, 12, 'local_g3_1')
// (16, 12, 'lutff_1/in_1')
// (16, 12, 'lutff_1/out')
// (16, 13, 'neigh_op_bot_1')
// (17, 11, 'neigh_op_tnl_1')
// (17, 12, 'local_g1_1')
// (17, 12, 'lutff_6/in_2')
// (17, 12, 'neigh_op_lft_1')
// (17, 13, 'local_g2_1')
// (17, 13, 'lutff_3/in_0')
// (17, 13, 'neigh_op_bnl_1')

reg n99 = 0;
// (15, 11, 'neigh_op_tnr_2')
// (15, 12, 'neigh_op_rgt_2')
// (15, 13, 'neigh_op_bnr_2')
// (16, 11, 'neigh_op_top_2')
// (16, 12, 'local_g1_2')
// (16, 12, 'lutff_2/in_1')
// (16, 12, 'lutff_2/out')
// (16, 13, 'neigh_op_bot_2')
// (17, 11, 'neigh_op_tnl_2')
// (17, 12, 'local_g1_2')
// (17, 12, 'lutff_6/in_3')
// (17, 12, 'neigh_op_lft_2')
// (17, 13, 'local_g3_2')
// (17, 13, 'lutff_0/in_1')
// (17, 13, 'neigh_op_bnl_2')

reg n100 = 0;
// (15, 11, 'neigh_op_tnr_3')
// (15, 12, 'neigh_op_rgt_3')
// (15, 13, 'neigh_op_bnr_3')
// (16, 11, 'neigh_op_top_3')
// (16, 12, 'local_g1_3')
// (16, 12, 'lutff_3/in_1')
// (16, 12, 'lutff_3/out')
// (16, 13, 'neigh_op_bot_3')
// (17, 11, 'neigh_op_tnl_3')
// (17, 12, 'local_g0_3')
// (17, 12, 'lutff_1/in_2')
// (17, 12, 'lutff_6/in_1')
// (17, 12, 'neigh_op_lft_3')
// (17, 13, 'neigh_op_bnl_3')

reg n101 = 0;
// (15, 11, 'neigh_op_tnr_4')
// (15, 12, 'neigh_op_rgt_4')
// (15, 13, 'neigh_op_bnr_4')
// (16, 11, 'neigh_op_top_4')
// (16, 12, 'local_g2_4')
// (16, 12, 'lutff_4/in_2')
// (16, 12, 'lutff_4/out')
// (16, 13, 'neigh_op_bot_4')
// (17, 11, 'neigh_op_tnl_4')
// (17, 12, 'local_g1_4')
// (17, 12, 'lutff_4/in_3')
// (17, 12, 'lutff_5/in_0')
// (17, 12, 'neigh_op_lft_4')
// (17, 13, 'neigh_op_bnl_4')

reg n102 = 0;
// (15, 11, 'neigh_op_tnr_5')
// (15, 12, 'neigh_op_rgt_5')
// (15, 13, 'neigh_op_bnr_5')
// (16, 11, 'neigh_op_top_5')
// (16, 12, 'local_g3_5')
// (16, 12, 'lutff_5/in_1')
// (16, 12, 'lutff_5/out')
// (16, 13, 'neigh_op_bot_5')
// (17, 11, 'neigh_op_tnl_5')
// (17, 12, 'local_g0_5')
// (17, 12, 'local_g1_5')
// (17, 12, 'lutff_0/in_3')
// (17, 12, 'lutff_5/in_3')
// (17, 12, 'neigh_op_lft_5')
// (17, 13, 'neigh_op_bnl_5')

reg n103 = 0;
// (15, 11, 'neigh_op_tnr_6')
// (15, 12, 'neigh_op_rgt_6')
// (15, 13, 'neigh_op_bnr_6')
// (16, 11, 'neigh_op_top_6')
// (16, 12, 'local_g3_6')
// (16, 12, 'lutff_6/in_1')
// (16, 12, 'lutff_6/out')
// (16, 13, 'neigh_op_bot_6')
// (17, 11, 'neigh_op_tnl_6')
// (17, 12, 'local_g0_6')
// (17, 12, 'lutff_5/in_1')
// (17, 12, 'lutff_7/in_1')
// (17, 12, 'neigh_op_lft_6')
// (17, 13, 'neigh_op_bnl_6')

reg n104 = 0;
// (15, 11, 'neigh_op_tnr_7')
// (15, 12, 'neigh_op_rgt_7')
// (15, 13, 'neigh_op_bnr_7')
// (16, 11, 'neigh_op_top_7')
// (16, 12, 'local_g3_7')
// (16, 12, 'lutff_7/in_1')
// (16, 12, 'lutff_7/out')
// (16, 13, 'neigh_op_bot_7')
// (17, 11, 'neigh_op_tnl_7')
// (17, 12, 'local_g0_7')
// (17, 12, 'lutff_5/in_2')
// (17, 12, 'neigh_op_lft_7')
// (17, 13, 'local_g2_7')
// (17, 13, 'lutff_5/in_2')
// (17, 13, 'neigh_op_bnl_7')

reg n105 = 0;
// (15, 11, 'sp4_r_v_b_43')
// (15, 12, 'sp4_r_v_b_30')
// (15, 13, 'sp4_r_v_b_19')
// (15, 14, 'sp4_r_v_b_6')
// (16, 10, 'sp4_h_r_0')
// (16, 10, 'sp4_v_t_43')
// (16, 11, 'local_g2_3')
// (16, 11, 'lutff_1/in_2')
// (16, 11, 'sp4_v_b_43')
// (16, 12, 'sp4_v_b_30')
// (16, 13, 'sp4_v_b_19')
// (16, 14, 'sp4_v_b_6')
// (17, 9, 'neigh_op_tnr_4')
// (17, 10, 'neigh_op_rgt_4')
// (17, 10, 'sp4_h_r_13')
// (17, 11, 'local_g1_4')
// (17, 11, 'lutff_3/in_2')
// (17, 11, 'neigh_op_bnr_4')
// (18, 9, 'neigh_op_top_4')
// (18, 10, 'local_g1_4')
// (18, 10, 'lutff_4/out')
// (18, 10, 'lutff_5/in_2')
// (18, 10, 'sp4_h_r_24')
// (18, 11, 'neigh_op_bot_4')
// (19, 9, 'neigh_op_tnl_4')
// (19, 10, 'neigh_op_lft_4')
// (19, 10, 'sp4_h_r_37')
// (19, 11, 'neigh_op_bnl_4')
// (20, 10, 'sp4_h_l_37')

reg n106 = 0;
// (15, 13, 'neigh_op_tnr_2')
// (15, 14, 'neigh_op_rgt_2')
// (15, 15, 'neigh_op_bnr_2')
// (16, 13, 'neigh_op_top_2')
// (16, 14, 'local_g2_2')
// (16, 14, 'lutff_2/in_2')
// (16, 14, 'lutff_2/out')
// (16, 14, 'lutff_5/in_3')
// (16, 15, 'neigh_op_bot_2')
// (17, 13, 'neigh_op_tnl_2')
// (17, 14, 'neigh_op_lft_2')
// (17, 15, 'neigh_op_bnl_2')

reg n107 = 0;
// (15, 13, 'neigh_op_tnr_3')
// (15, 14, 'neigh_op_rgt_3')
// (15, 15, 'neigh_op_bnr_3')
// (16, 13, 'neigh_op_top_3')
// (16, 14, 'local_g3_3')
// (16, 14, 'lutff_0/in_2')
// (16, 14, 'lutff_3/in_3')
// (16, 14, 'lutff_3/out')
// (16, 14, 'lutff_5/in_1')
// (16, 15, 'local_g0_3')
// (16, 15, 'lutff_2/in_3')
// (16, 15, 'neigh_op_bot_3')
// (17, 13, 'neigh_op_tnl_3')
// (17, 14, 'neigh_op_lft_3')
// (17, 15, 'neigh_op_bnl_3')

wire n108;
// (15, 13, 'neigh_op_tnr_4')
// (15, 14, 'neigh_op_rgt_4')
// (15, 15, 'neigh_op_bnr_4')
// (16, 13, 'neigh_op_top_4')
// (16, 14, 'local_g0_4')
// (16, 14, 'local_g1_4')
// (16, 14, 'lutff_4/out')
// (16, 14, 'lutff_5/in_0')
// (16, 14, 'lutff_global/s_r')
// (16, 15, 'local_g0_4')
// (16, 15, 'lutff_2/in_2')
// (16, 15, 'lutff_global/s_r')
// (16, 15, 'neigh_op_bot_4')
// (17, 13, 'neigh_op_tnl_4')
// (17, 14, 'neigh_op_lft_4')
// (17, 15, 'neigh_op_bnl_4')

wire n109;
// (15, 14, 'neigh_op_tnr_2')
// (15, 15, 'neigh_op_rgt_2')
// (15, 16, 'neigh_op_bnr_2')
// (16, 14, 'neigh_op_top_2')
// (16, 15, 'local_g2_2')
// (16, 15, 'lutff_2/out')
// (16, 15, 'lutff_global/cen')
// (16, 16, 'neigh_op_bot_2')
// (17, 14, 'neigh_op_tnl_2')
// (17, 15, 'neigh_op_lft_2')
// (17, 16, 'neigh_op_bnl_2')

reg n110 = 0;
// (15, 14, 'neigh_op_tnr_3')
// (15, 15, 'neigh_op_rgt_3')
// (15, 16, 'neigh_op_bnr_3')
// (16, 14, 'local_g0_3')
// (16, 14, 'lutff_1/in_2')
// (16, 14, 'lutff_5/in_2')
// (16, 14, 'neigh_op_top_3')
// (16, 15, 'local_g1_3')
// (16, 15, 'lutff_3/in_3')
// (16, 15, 'lutff_3/out')
// (16, 16, 'neigh_op_bot_3')
// (17, 14, 'neigh_op_tnl_3')
// (17, 15, 'neigh_op_lft_3')
// (17, 16, 'neigh_op_bnl_3')

wire n111;
// (16, 9, 'neigh_op_tnr_2')
// (16, 10, 'neigh_op_rgt_2')
// (16, 11, 'neigh_op_bnr_2')
// (17, 9, 'neigh_op_top_2')
// (17, 10, 'lutff_2/out')
// (17, 11, 'neigh_op_bot_2')
// (18, 9, 'neigh_op_tnl_2')
// (18, 10, 'neigh_op_lft_2')
// (18, 11, 'local_g2_2')
// (18, 11, 'lutff_2/in_2')
// (18, 11, 'neigh_op_bnl_2')

wire n112;
// (16, 9, 'neigh_op_tnr_3')
// (16, 10, 'neigh_op_rgt_3')
// (16, 11, 'neigh_op_bnr_3')
// (17, 9, 'neigh_op_top_3')
// (17, 10, 'lutff_3/out')
// (17, 11, 'neigh_op_bot_3')
// (18, 9, 'neigh_op_tnl_3')
// (18, 10, 'neigh_op_lft_3')
// (18, 11, 'local_g3_3')
// (18, 11, 'lutff_4/in_2')
// (18, 11, 'neigh_op_bnl_3')

wire n113;
// (16, 10, 'neigh_op_tnr_0')
// (16, 11, 'neigh_op_rgt_0')
// (16, 12, 'neigh_op_bnr_0')
// (17, 10, 'neigh_op_top_0')
// (17, 11, 'lutff_0/out')
// (17, 12, 'neigh_op_bot_0')
// (18, 10, 'neigh_op_tnl_0')
// (18, 11, 'local_g1_0')
// (18, 11, 'lutff_6/in_1')
// (18, 11, 'neigh_op_lft_0')
// (18, 12, 'neigh_op_bnl_0')

wire n114;
// (16, 10, 'neigh_op_tnr_1')
// (16, 11, 'neigh_op_rgt_1')
// (16, 12, 'neigh_op_bnr_1')
// (17, 10, 'neigh_op_top_1')
// (17, 11, 'lutff_1/out')
// (17, 12, 'neigh_op_bot_1')
// (18, 10, 'neigh_op_tnl_1')
// (18, 11, 'local_g1_1')
// (18, 11, 'lutff_5/in_1')
// (18, 11, 'neigh_op_lft_1')
// (18, 12, 'neigh_op_bnl_1')

wire n115;
// (16, 10, 'neigh_op_tnr_2')
// (16, 11, 'neigh_op_rgt_2')
// (16, 12, 'neigh_op_bnr_2')
// (17, 10, 'neigh_op_top_2')
// (17, 11, 'lutff_2/out')
// (17, 12, 'local_g0_2')
// (17, 12, 'lutff_2/in_0')
// (17, 12, 'neigh_op_bot_2')
// (18, 10, 'neigh_op_tnl_2')
// (18, 11, 'neigh_op_lft_2')
// (18, 12, 'neigh_op_bnl_2')

wire n116;
// (16, 10, 'neigh_op_tnr_3')
// (16, 11, 'neigh_op_rgt_3')
// (16, 12, 'neigh_op_bnr_3')
// (17, 10, 'neigh_op_top_3')
// (17, 11, 'lutff_3/out')
// (17, 12, 'local_g1_3')
// (17, 12, 'lutff_2/in_2')
// (17, 12, 'neigh_op_bot_3')
// (18, 10, 'neigh_op_tnl_3')
// (18, 11, 'neigh_op_lft_3')
// (18, 12, 'neigh_op_bnl_3')

wire n117;
// (16, 10, 'neigh_op_tnr_4')
// (16, 11, 'neigh_op_rgt_4')
// (16, 12, 'neigh_op_bnr_4')
// (17, 10, 'neigh_op_top_4')
// (17, 11, 'lutff_4/out')
// (17, 12, 'neigh_op_bot_4')
// (18, 10, 'neigh_op_tnl_4')
// (18, 11, 'local_g0_4')
// (18, 11, 'lutff_3/in_1')
// (18, 11, 'neigh_op_lft_4')
// (18, 12, 'neigh_op_bnl_4')

wire n118;
// (16, 10, 'neigh_op_tnr_5')
// (16, 11, 'neigh_op_rgt_5')
// (16, 12, 'neigh_op_bnr_5')
// (17, 10, 'neigh_op_top_5')
// (17, 11, 'lutff_5/out')
// (17, 12, 'neigh_op_bot_5')
// (18, 10, 'neigh_op_tnl_5')
// (18, 11, 'local_g1_5')
// (18, 11, 'lutff_7/in_1')
// (18, 11, 'neigh_op_lft_5')
// (18, 12, 'neigh_op_bnl_5')

reg n119 = 0;
// (16, 10, 'neigh_op_tnr_7')
// (16, 11, 'local_g3_7')
// (16, 11, 'lutff_0/in_2')
// (16, 11, 'neigh_op_rgt_7')
// (16, 12, 'neigh_op_bnr_7')
// (17, 10, 'neigh_op_top_7')
// (17, 11, 'local_g1_7')
// (17, 11, 'lutff_3/in_3')
// (17, 11, 'lutff_7/in_3')
// (17, 11, 'lutff_7/out')
// (17, 12, 'neigh_op_bot_7')
// (18, 10, 'local_g2_7')
// (18, 10, 'local_g3_7')
// (18, 10, 'lutff_0/in_2')
// (18, 10, 'lutff_7/in_2')
// (18, 10, 'neigh_op_tnl_7')
// (18, 11, 'neigh_op_lft_7')
// (18, 12, 'neigh_op_bnl_7')

wire n120;
// (16, 10, 'sp4_r_v_b_42')
// (16, 11, 'sp4_r_v_b_31')
// (16, 12, 'sp4_r_v_b_18')
// (16, 13, 'sp4_r_v_b_7')
// (16, 14, 'sp4_r_v_b_41')
// (16, 15, 'sp4_r_v_b_28')
// (16, 16, 'sp4_r_v_b_17')
// (16, 17, 'sp4_r_v_b_4')
// (16, 18, 'sp4_r_v_b_45')
// (16, 19, 'sp4_r_v_b_32')
// (16, 20, 'neigh_op_tnr_4')
// (16, 20, 'sp4_r_v_b_21')
// (16, 21, 'neigh_op_rgt_4')
// (16, 21, 'sp4_r_v_b_8')
// (16, 22, 'neigh_op_bnr_4')
// (17, 9, 'sp4_v_t_42')
// (17, 10, 'sp4_v_b_42')
// (17, 11, 'local_g2_7')
// (17, 11, 'lutff_6/in_1')
// (17, 11, 'sp4_v_b_31')
// (17, 12, 'sp4_v_b_18')
// (17, 13, 'sp4_v_b_7')
// (17, 13, 'sp4_v_t_41')
// (17, 14, 'sp4_v_b_41')
// (17, 15, 'sp4_v_b_28')
// (17, 16, 'sp4_v_b_17')
// (17, 17, 'sp4_v_b_4')
// (17, 17, 'sp4_v_t_45')
// (17, 18, 'sp4_v_b_45')
// (17, 19, 'sp4_v_b_32')
// (17, 20, 'neigh_op_top_4')
// (17, 20, 'sp4_v_b_21')
// (17, 21, 'lutff_4/out')
// (17, 21, 'sp4_v_b_8')
// (17, 22, 'neigh_op_bot_4')
// (18, 20, 'neigh_op_tnl_4')
// (18, 21, 'neigh_op_lft_4')
// (18, 22, 'neigh_op_bnl_4')

wire n121;
// (16, 11, 'local_g3_3')
// (16, 11, 'lutff_global/cen')
// (16, 11, 'neigh_op_tnr_3')
// (16, 12, 'local_g3_3')
// (16, 12, 'lutff_global/cen')
// (16, 12, 'neigh_op_rgt_3')
// (16, 13, 'neigh_op_bnr_3')
// (17, 11, 'local_g1_3')
// (17, 11, 'lutff_global/cen')
// (17, 11, 'neigh_op_top_3')
// (17, 12, 'lutff_3/out')
// (17, 13, 'neigh_op_bot_3')
// (18, 11, 'neigh_op_tnl_3')
// (18, 12, 'neigh_op_lft_3')
// (18, 13, 'neigh_op_bnl_3')

wire n122;
// (16, 11, 'lutff_1/cout')
// (16, 11, 'lutff_2/in_3')

wire n123;
// (16, 11, 'lutff_2/cout')
// (16, 11, 'lutff_3/in_3')

wire n124;
// (16, 11, 'lutff_3/cout')
// (16, 11, 'lutff_4/in_3')

wire n125;
// (16, 11, 'lutff_4/cout')
// (16, 11, 'lutff_5/in_3')

wire n126;
// (16, 11, 'lutff_5/cout')
// (16, 11, 'lutff_6/in_3')

wire n127;
// (16, 11, 'lutff_6/cout')
// (16, 11, 'lutff_7/in_3')

wire n128;
// (16, 11, 'lutff_7/cout')
// (16, 12, 'carry_in')
// (16, 12, 'carry_in_mux')
// (16, 12, 'lutff_0/in_3')

wire n129;
// (16, 11, 'neigh_op_tnr_0')
// (16, 12, 'neigh_op_rgt_0')
// (16, 13, 'neigh_op_bnr_0')
// (17, 11, 'neigh_op_top_0')
// (17, 12, 'lutff_0/out')
// (17, 13, 'neigh_op_bot_0')
// (18, 11, 'neigh_op_tnl_0')
// (18, 12, 'local_g1_0')
// (18, 12, 'lutff_5/in_2')
// (18, 12, 'neigh_op_lft_0')
// (18, 13, 'neigh_op_bnl_0')

wire n130;
// (16, 11, 'neigh_op_tnr_1')
// (16, 12, 'neigh_op_rgt_1')
// (16, 13, 'neigh_op_bnr_1')
// (17, 11, 'neigh_op_top_1')
// (17, 12, 'lutff_1/out')
// (17, 13, 'neigh_op_bot_1')
// (18, 11, 'neigh_op_tnl_1')
// (18, 12, 'local_g1_1')
// (18, 12, 'lutff_3/in_1')
// (18, 12, 'neigh_op_lft_1')
// (18, 13, 'neigh_op_bnl_1')

wire n131;
// (16, 11, 'neigh_op_tnr_2')
// (16, 12, 'neigh_op_rgt_2')
// (16, 13, 'neigh_op_bnr_2')
// (17, 11, 'local_g1_2')
// (17, 11, 'lutff_6/in_3')
// (17, 11, 'neigh_op_top_2')
// (17, 12, 'lutff_2/out')
// (17, 13, 'neigh_op_bot_2')
// (18, 11, 'neigh_op_tnl_2')
// (18, 12, 'neigh_op_lft_2')
// (18, 13, 'neigh_op_bnl_2')

wire n132;
// (16, 11, 'neigh_op_tnr_4')
// (16, 12, 'neigh_op_rgt_4')
// (16, 13, 'neigh_op_bnr_4')
// (17, 11, 'neigh_op_top_4')
// (17, 12, 'lutff_4/out')
// (17, 13, 'neigh_op_bot_4')
// (18, 11, 'neigh_op_tnl_4')
// (18, 12, 'local_g0_4')
// (18, 12, 'lutff_4/in_2')
// (18, 12, 'neigh_op_lft_4')
// (18, 13, 'neigh_op_bnl_4')

wire n133;
// (16, 11, 'neigh_op_tnr_5')
// (16, 12, 'neigh_op_rgt_5')
// (16, 13, 'neigh_op_bnr_5')
// (17, 11, 'neigh_op_top_5')
// (17, 12, 'local_g2_5')
// (17, 12, 'lutff_2/in_1')
// (17, 12, 'lutff_5/out')
// (17, 13, 'neigh_op_bot_5')
// (18, 11, 'neigh_op_tnl_5')
// (18, 12, 'neigh_op_lft_5')
// (18, 13, 'neigh_op_bnl_5')

wire n134;
// (16, 11, 'neigh_op_tnr_6')
// (16, 12, 'neigh_op_rgt_6')
// (16, 13, 'neigh_op_bnr_6')
// (17, 11, 'neigh_op_top_6')
// (17, 12, 'local_g3_6')
// (17, 12, 'lutff_2/in_3')
// (17, 12, 'lutff_6/out')
// (17, 13, 'neigh_op_bot_6')
// (18, 11, 'neigh_op_tnl_6')
// (18, 12, 'neigh_op_lft_6')
// (18, 13, 'neigh_op_bnl_6')

wire n135;
// (16, 11, 'neigh_op_tnr_7')
// (16, 12, 'neigh_op_rgt_7')
// (16, 13, 'neigh_op_bnr_7')
// (17, 11, 'neigh_op_top_7')
// (17, 12, 'lutff_7/out')
// (17, 13, 'neigh_op_bot_7')
// (18, 11, 'neigh_op_tnl_7')
// (18, 12, 'local_g0_7')
// (18, 12, 'lutff_6/in_1')
// (18, 12, 'neigh_op_lft_7')
// (18, 13, 'neigh_op_bnl_7')

wire n136;
// (16, 12, 'lutff_0/cout')
// (16, 12, 'lutff_1/in_3')

wire n137;
// (16, 12, 'lutff_1/cout')
// (16, 12, 'lutff_2/in_3')

wire n138;
// (16, 12, 'lutff_2/cout')
// (16, 12, 'lutff_3/in_3')

wire n139;
// (16, 12, 'lutff_3/cout')
// (16, 12, 'lutff_4/in_3')

wire n140;
// (16, 12, 'lutff_4/cout')
// (16, 12, 'lutff_5/in_3')

wire n141;
// (16, 12, 'lutff_5/cout')
// (16, 12, 'lutff_6/in_3')

wire n142;
// (16, 12, 'lutff_6/cout')
// (16, 12, 'lutff_7/in_3')

wire n143;
// (16, 12, 'neigh_op_tnr_0')
// (16, 13, 'neigh_op_rgt_0')
// (16, 14, 'neigh_op_bnr_0')
// (17, 12, 'neigh_op_top_0')
// (17, 13, 'lutff_0/out')
// (17, 14, 'neigh_op_bot_0')
// (18, 12, 'local_g2_0')
// (18, 12, 'lutff_2/in_2')
// (18, 12, 'neigh_op_tnl_0')
// (18, 13, 'neigh_op_lft_0')
// (18, 14, 'neigh_op_bnl_0')

wire n144;
// (16, 12, 'neigh_op_tnr_3')
// (16, 13, 'neigh_op_rgt_3')
// (16, 14, 'neigh_op_bnr_3')
// (17, 12, 'neigh_op_top_3')
// (17, 13, 'lutff_3/out')
// (17, 14, 'neigh_op_bot_3')
// (18, 12, 'local_g2_3')
// (18, 12, 'lutff_1/in_2')
// (18, 12, 'neigh_op_tnl_3')
// (18, 13, 'neigh_op_lft_3')
// (18, 14, 'neigh_op_bnl_3')

wire n145;
// (16, 12, 'neigh_op_tnr_5')
// (16, 13, 'neigh_op_rgt_5')
// (16, 14, 'neigh_op_bnr_5')
// (17, 12, 'neigh_op_top_5')
// (17, 13, 'lutff_5/out')
// (17, 14, 'neigh_op_bot_5')
// (18, 12, 'local_g2_5')
// (18, 12, 'lutff_7/in_2')
// (18, 12, 'neigh_op_tnl_5')
// (18, 13, 'neigh_op_lft_5')
// (18, 14, 'neigh_op_bnl_5')

wire n146;
// (16, 12, 'neigh_op_tnr_7')
// (16, 13, 'neigh_op_rgt_7')
// (16, 14, 'neigh_op_bnr_7')
// (17, 12, 'neigh_op_top_7')
// (17, 13, 'lutff_7/out')
// (17, 14, 'neigh_op_bot_7')
// (18, 12, 'local_g3_7')
// (18, 12, 'lutff_0/in_2')
// (18, 12, 'neigh_op_tnl_7')
// (18, 13, 'neigh_op_lft_7')
// (18, 14, 'neigh_op_bnl_7')

wire n147;
// (16, 14, 'lutff_1/cout')
// (16, 14, 'lutff_2/in_3')

wire io_29_0_0;
// (17, 5, 'sp12_h_r_0')
// (17, 5, 'sp12_v_t_23')
// (17, 6, 'sp12_v_b_23')
// (17, 7, 'sp12_v_b_20')
// (17, 8, 'sp12_v_b_19')
// (17, 9, 'sp12_v_b_16')
// (17, 10, 'sp12_v_b_15')
// (17, 11, 'local_g2_4')
// (17, 11, 'lutff_6/in_2')
// (17, 11, 'sp12_v_b_12')
// (17, 12, 'sp12_v_b_11')
// (17, 13, 'sp12_v_b_8')
// (17, 14, 'sp12_v_b_7')
// (17, 15, 'sp12_v_b_4')
// (17, 16, 'sp12_v_b_3')
// (17, 17, 'sp12_v_b_0')
// (18, 5, 'sp12_h_r_3')
// (19, 5, 'sp12_h_r_4')
// (20, 5, 'sp12_h_r_7')
// (21, 5, 'sp12_h_r_8')
// (22, 5, 'sp12_h_r_11')
// (23, 5, 'sp12_h_r_12')
// (24, 5, 'sp12_h_r_15')
// (25, 5, 'sp12_h_r_16')
// (26, 5, 'sp12_h_r_19')
// (27, 5, 'sp12_h_r_20')
// (28, 1, 'neigh_op_bnr_0')
// (28, 1, 'neigh_op_bnr_4')
// (28, 5, 'sp12_h_r_23')
// (29, 0, 'io_0/D_IN_0')
// (29, 0, 'io_0/PAD')
// (29, 0, 'span12_vert_8')
// (29, 1, 'neigh_op_bot_0')
// (29, 1, 'neigh_op_bot_4')
// (29, 1, 'sp12_v_b_8')
// (29, 2, 'sp12_v_b_7')
// (29, 3, 'sp12_v_b_4')
// (29, 4, 'sp12_v_b_3')
// (29, 5, 'sp12_h_l_23')
// (29, 5, 'sp12_v_b_0')
// (30, 1, 'neigh_op_bnl_0')
// (30, 1, 'neigh_op_bnl_4')

wire n149;
// (17, 9, 'neigh_op_tnr_0')
// (17, 10, 'neigh_op_rgt_0')
// (17, 11, 'neigh_op_bnr_0')
// (18, 9, 'neigh_op_top_0')
// (18, 10, 'lutff_0/out')
// (18, 11, 'local_g0_0')
// (18, 11, 'lutff_0/in_2')
// (18, 11, 'neigh_op_bot_0')
// (19, 9, 'neigh_op_tnl_0')
// (19, 10, 'neigh_op_lft_0')
// (19, 11, 'neigh_op_bnl_0')

wire n150;
// (17, 9, 'neigh_op_tnr_2')
// (17, 10, 'neigh_op_rgt_2')
// (17, 11, 'neigh_op_bnr_2')
// (18, 9, 'neigh_op_top_2')
// (18, 10, 'local_g0_2')
// (18, 10, 'lutff_2/out')
// (18, 10, 'lutff_global/cen')
// (18, 11, 'neigh_op_bot_2')
// (19, 9, 'neigh_op_tnl_2')
// (19, 10, 'neigh_op_lft_2')
// (19, 11, 'neigh_op_bnl_2')

wire n151;
// (17, 9, 'neigh_op_tnr_5')
// (17, 10, 'neigh_op_rgt_5')
// (17, 11, 'neigh_op_bnr_5')
// (18, 9, 'neigh_op_top_5')
// (18, 10, 'local_g1_5')
// (18, 10, 'lutff_4/in_0')
// (18, 10, 'lutff_5/out')
// (18, 11, 'local_g0_5')
// (18, 11, 'lutff_1/in_2')
// (18, 11, 'neigh_op_bot_5')
// (19, 9, 'neigh_op_tnl_5')
// (19, 10, 'neigh_op_lft_5')
// (19, 11, 'neigh_op_bnl_5')

wire n152;
// (17, 9, 'neigh_op_tnr_7')
// (17, 10, 'neigh_op_rgt_7')
// (17, 11, 'neigh_op_bnr_7')
// (18, 9, 'neigh_op_top_7')
// (18, 10, 'local_g0_7')
// (18, 10, 'lutff_2/in_1')
// (18, 10, 'lutff_7/out')
// (18, 11, 'neigh_op_bot_7')
// (19, 9, 'neigh_op_tnl_7')
// (19, 10, 'neigh_op_lft_7')
// (19, 11, 'neigh_op_bnl_7')

wire n153;
// (17, 10, 'sp4_r_v_b_36')
// (17, 11, 'local_g1_1')
// (17, 11, 'lutff_6/in_0')
// (17, 11, 'sp4_r_v_b_25')
// (17, 12, 'sp4_r_v_b_12')
// (17, 13, 'sp4_r_v_b_1')
// (18, 9, 'sp4_v_t_36')
// (18, 10, 'sp4_v_b_36')
// (18, 11, 'sp4_v_b_25')
// (18, 12, 'sp4_v_b_12')
// (18, 13, 'sp4_h_r_8')
// (18, 13, 'sp4_v_b_1')
// (19, 13, 'sp4_h_r_21')
// (20, 13, 'sp4_h_r_32')
// (21, 13, 'sp4_h_r_45')
// (21, 14, 'sp4_r_v_b_45')
// (21, 15, 'sp4_r_v_b_32')
// (21, 16, 'sp4_r_v_b_21')
// (21, 17, 'sp4_r_v_b_8')
// (21, 18, 'sp4_r_v_b_45')
// (21, 19, 'sp4_r_v_b_32')
// (21, 20, 'neigh_op_tnr_4')
// (21, 20, 'sp4_r_v_b_21')
// (21, 21, 'neigh_op_rgt_4')
// (21, 21, 'sp4_r_v_b_8')
// (21, 22, 'neigh_op_bnr_4')
// (22, 13, 'sp4_h_l_45')
// (22, 13, 'sp4_v_t_45')
// (22, 14, 'sp4_v_b_45')
// (22, 15, 'sp4_v_b_32')
// (22, 16, 'sp4_v_b_21')
// (22, 17, 'sp4_v_b_8')
// (22, 17, 'sp4_v_t_45')
// (22, 18, 'sp4_v_b_45')
// (22, 19, 'sp4_v_b_32')
// (22, 20, 'neigh_op_top_4')
// (22, 20, 'sp4_v_b_21')
// (22, 21, 'lutff_4/out')
// (22, 21, 'sp4_v_b_8')
// (22, 22, 'neigh_op_bot_4')
// (23, 20, 'neigh_op_tnl_4')
// (23, 21, 'neigh_op_lft_4')
// (23, 22, 'neigh_op_bnl_4')

wire n154;
// (17, 10, 'sp4_r_v_b_37')
// (17, 11, 'sp4_r_v_b_24')
// (17, 12, 'local_g2_0')
// (17, 12, 'lutff_3/in_1')
// (17, 12, 'neigh_op_tnr_0')
// (17, 12, 'sp4_r_v_b_13')
// (17, 13, 'neigh_op_rgt_0')
// (17, 13, 'sp4_r_v_b_0')
// (17, 14, 'neigh_op_bnr_0')
// (18, 9, 'sp4_v_t_37')
// (18, 10, 'local_g3_5')
// (18, 10, 'lutff_7/in_3')
// (18, 10, 'sp4_v_b_37')
// (18, 11, 'sp4_v_b_24')
// (18, 12, 'neigh_op_top_0')
// (18, 12, 'sp4_v_b_13')
// (18, 13, 'lutff_0/out')
// (18, 13, 'sp4_v_b_0')
// (18, 14, 'neigh_op_bot_0')
// (19, 12, 'local_g2_0')
// (19, 12, 'lutff_5/in_3')
// (19, 12, 'neigh_op_tnl_0')
// (19, 13, 'neigh_op_lft_0')
// (19, 14, 'neigh_op_bnl_0')

wire n155;
// (17, 21, 'local_g0_0')
// (17, 21, 'lutff_4/in_0')
// (17, 21, 'sp12_h_r_0')
// (18, 21, 'sp12_h_r_3')
// (19, 21, 'sp12_h_r_4')
// (20, 20, 'neigh_op_tnr_0')
// (20, 21, 'neigh_op_rgt_0')
// (20, 21, 'sp12_h_r_7')
// (20, 22, 'neigh_op_bnr_0')
// (21, 20, 'neigh_op_top_0')
// (21, 21, 'lutff_0/out')
// (21, 21, 'sp12_h_r_8')
// (21, 22, 'neigh_op_bot_0')
// (22, 20, 'neigh_op_tnl_0')
// (22, 21, 'neigh_op_lft_0')
// (22, 21, 'sp12_h_r_11')
// (22, 22, 'neigh_op_bnl_0')
// (23, 21, 'sp12_h_r_12')
// (24, 21, 'sp12_h_r_15')
// (25, 21, 'sp12_h_r_16')
// (26, 21, 'sp12_h_r_19')
// (27, 21, 'sp12_h_r_20')
// (28, 21, 'sp12_h_r_23')
// (29, 21, 'sp12_h_l_23')

wire n156;
// (18, 11, 'lutff_7/cout')
// (18, 12, 'carry_in')
// (18, 12, 'carry_in_mux')

wire n157;
// (18, 11, 'neigh_op_tnr_5')
// (18, 12, 'neigh_op_rgt_5')
// (18, 12, 'sp12_h_r_1')
// (18, 13, 'neigh_op_bnr_5')
// (19, 11, 'neigh_op_top_5')
// (19, 12, 'lutff_5/out')
// (19, 12, 'sp12_h_r_2')
// (19, 13, 'neigh_op_bot_5')
// (20, 11, 'neigh_op_tnl_5')
// (20, 12, 'neigh_op_lft_5')
// (20, 12, 'sp12_h_r_5')
// (20, 13, 'neigh_op_bnl_5')
// (21, 12, 'sp12_h_r_6')
// (22, 12, 'sp12_h_r_9')
// (23, 12, 'sp12_h_r_10')
// (24, 12, 'sp12_h_r_13')
// (25, 12, 'sp12_h_r_14')
// (26, 12, 'sp12_h_r_17')
// (27, 12, 'sp12_h_r_18')
// (28, 12, 'sp12_h_r_21')
// (29, 12, 'sp12_h_r_22')
// (30, 0, 'span12_vert_22')
// (30, 1, 'local_g3_6')
// (30, 1, 'lutff_6/in_1')
// (30, 1, 'sp12_v_b_22')
// (30, 2, 'sp12_v_b_21')
// (30, 3, 'sp12_v_b_18')
// (30, 4, 'sp12_v_b_17')
// (30, 5, 'sp12_v_b_14')
// (30, 6, 'sp12_v_b_13')
// (30, 7, 'sp12_v_b_10')
// (30, 8, 'sp12_v_b_9')
// (30, 9, 'sp12_v_b_6')
// (30, 10, 'sp12_v_b_5')
// (30, 11, 'sp12_v_b_2')
// (30, 12, 'sp12_h_l_22')
// (30, 12, 'sp12_v_b_1')

wire n158;
// (18, 12, 'lutff_7/cout')
// (18, 13, 'carry_in')
// (18, 13, 'carry_in_mux')
// (18, 13, 'lutff_0/in_3')

wire n159;
// (19, 18, 'neigh_op_tnr_5')
// (19, 19, 'neigh_op_rgt_5')
// (19, 20, 'neigh_op_bnr_5')
// (20, 18, 'neigh_op_top_5')
// (20, 19, 'lutff_5/out')
// (20, 19, 'sp4_h_r_10')
// (20, 20, 'neigh_op_bot_5')
// (21, 18, 'neigh_op_tnl_5')
// (21, 19, 'local_g1_5')
// (21, 19, 'lutff_7/in_1')
// (21, 19, 'neigh_op_lft_5')
// (21, 19, 'sp4_h_r_23')
// (21, 20, 'neigh_op_bnl_5')
// (22, 19, 'local_g3_2')
// (22, 19, 'lutff_7/in_2')
// (22, 19, 'sp4_h_r_34')
// (23, 19, 'sp4_h_r_47')
// (24, 19, 'sp4_h_l_47')

wire n160;
// (19, 18, 'neigh_op_tnr_6')
// (19, 19, 'neigh_op_rgt_6')
// (19, 19, 'sp4_h_r_1')
// (19, 20, 'neigh_op_bnr_6')
// (20, 18, 'neigh_op_top_6')
// (20, 19, 'lutff_6/out')
// (20, 19, 'sp4_h_r_12')
// (20, 20, 'neigh_op_bot_6')
// (21, 18, 'neigh_op_tnl_6')
// (21, 19, 'local_g1_6')
// (21, 19, 'lutff_4/in_1')
// (21, 19, 'neigh_op_lft_6')
// (21, 19, 'sp4_h_r_25')
// (21, 20, 'neigh_op_bnl_6')
// (22, 19, 'local_g2_4')
// (22, 19, 'lutff_4/in_2')
// (22, 19, 'sp4_h_r_36')
// (23, 19, 'sp4_h_l_36')

wire n161;
// (19, 18, 'neigh_op_tnr_7')
// (19, 19, 'neigh_op_rgt_7')
// (19, 19, 'sp4_h_r_3')
// (19, 20, 'neigh_op_bnr_7')
// (20, 18, 'neigh_op_top_7')
// (20, 19, 'lutff_7/out')
// (20, 19, 'sp4_h_r_14')
// (20, 20, 'neigh_op_bot_7')
// (21, 18, 'neigh_op_tnl_7')
// (21, 19, 'local_g1_7')
// (21, 19, 'lutff_5/in_1')
// (21, 19, 'neigh_op_lft_7')
// (21, 19, 'sp4_h_r_27')
// (21, 20, 'neigh_op_bnl_7')
// (22, 19, 'local_g2_6')
// (22, 19, 'lutff_5/in_1')
// (22, 19, 'sp4_h_r_38')
// (23, 19, 'sp4_h_l_38')

wire n162;
// (19, 19, 'neigh_op_tnr_2')
// (19, 20, 'neigh_op_rgt_2')
// (19, 21, 'neigh_op_bnr_2')
// (20, 19, 'neigh_op_top_2')
// (20, 20, 'lutff_2/out')
// (20, 20, 'sp4_h_r_4')
// (20, 21, 'neigh_op_bot_2')
// (21, 19, 'neigh_op_tnl_2')
// (21, 20, 'local_g0_2')
// (21, 20, 'lutff_1/in_1')
// (21, 20, 'neigh_op_lft_2')
// (21, 20, 'sp4_h_r_17')
// (21, 21, 'neigh_op_bnl_2')
// (22, 20, 'local_g2_4')
// (22, 20, 'lutff_1/in_1')
// (22, 20, 'sp4_h_r_28')
// (23, 20, 'sp4_h_r_41')
// (24, 20, 'sp4_h_l_41')

wire n163;
// (20, 17, 'neigh_op_tnr_3')
// (20, 18, 'neigh_op_rgt_3')
// (20, 19, 'neigh_op_bnr_3')
// (21, 17, 'neigh_op_top_3')
// (21, 18, 'lutff_3/out')
// (21, 19, 'local_g1_3')
// (21, 19, 'lutff_1/in_1')
// (21, 19, 'neigh_op_bot_3')
// (22, 17, 'neigh_op_tnl_3')
// (22, 18, 'neigh_op_lft_3')
// (22, 19, 'local_g3_3')
// (22, 19, 'lutff_1/in_1')
// (22, 19, 'neigh_op_bnl_3')

wire n164;
// (20, 18, 'sp4_r_v_b_38')
// (20, 19, 'sp4_r_v_b_27')
// (20, 20, 'sp4_r_v_b_14')
// (20, 21, 'sp4_r_v_b_3')
// (21, 17, 'sp4_v_t_38')
// (21, 18, 'sp4_v_b_38')
// (21, 19, 'sp4_v_b_27')
// (21, 20, 'local_g1_6')
// (21, 20, 'lutff_7/in_2')
// (21, 20, 'sp4_v_b_14')
// (21, 21, 'sp4_h_r_3')
// (21, 21, 'sp4_v_b_3')
// (22, 18, 'sp4_r_v_b_41')
// (22, 19, 'sp4_r_v_b_28')
// (22, 20, 'local_g3_1')
// (22, 20, 'lutff_7/in_1')
// (22, 20, 'sp4_r_v_b_17')
// (22, 21, 'sp4_h_r_14')
// (22, 21, 'sp4_r_v_b_4')
// (23, 17, 'sp4_v_t_41')
// (23, 18, 'sp4_v_b_41')
// (23, 19, 'sp4_v_b_28')
// (23, 20, 'neigh_op_tnr_3')
// (23, 20, 'sp4_v_b_17')
// (23, 21, 'neigh_op_rgt_3')
// (23, 21, 'sp4_h_r_11')
// (23, 21, 'sp4_h_r_27')
// (23, 21, 'sp4_v_b_4')
// (23, 22, 'neigh_op_bnr_3')
// (24, 20, 'neigh_op_top_3')
// (24, 21, 'lutff_3/out')
// (24, 21, 'sp4_h_r_22')
// (24, 21, 'sp4_h_r_38')
// (24, 22, 'neigh_op_bot_3')
// (25, 20, 'neigh_op_tnl_3')
// (25, 21, 'neigh_op_lft_3')
// (25, 21, 'sp4_h_l_38')
// (25, 21, 'sp4_h_r_35')
// (25, 22, 'neigh_op_bnl_3')
// (26, 21, 'sp4_h_r_46')
// (27, 21, 'sp4_h_l_46')

wire n165;
// (20, 20, 'sp4_h_r_0')
// (21, 20, 'local_g0_5')
// (21, 20, 'lutff_4/in_1')
// (21, 20, 'sp4_h_r_13')
// (22, 17, 'sp4_r_v_b_44')
// (22, 18, 'sp4_r_v_b_33')
// (22, 19, 'sp4_r_v_b_20')
// (22, 20, 'local_g2_1')
// (22, 20, 'lutff_4/in_1')
// (22, 20, 'sp4_h_r_24')
// (22, 20, 'sp4_r_v_b_9')
// (23, 16, 'sp4_v_t_44')
// (23, 17, 'sp4_v_b_44')
// (23, 18, 'sp4_v_b_33')
// (23, 19, 'sp4_v_b_20')
// (23, 20, 'sp4_h_r_37')
// (23, 20, 'sp4_h_r_9')
// (23, 20, 'sp4_v_b_9')
// (24, 20, 'sp4_h_l_37')
// (24, 20, 'sp4_h_r_20')
// (24, 20, 'sp4_h_r_4')
// (25, 19, 'neigh_op_tnr_6')
// (25, 20, 'neigh_op_rgt_6')
// (25, 20, 'sp4_h_r_17')
// (25, 20, 'sp4_h_r_33')
// (25, 21, 'neigh_op_bnr_6')
// (26, 19, 'neigh_op_top_6')
// (26, 20, 'lutff_6/out')
// (26, 20, 'sp4_h_r_28')
// (26, 20, 'sp4_h_r_44')
// (26, 21, 'neigh_op_bot_6')
// (27, 19, 'neigh_op_tnl_6')
// (27, 20, 'neigh_op_lft_6')
// (27, 20, 'sp4_h_l_44')
// (27, 20, 'sp4_h_r_41')
// (27, 21, 'neigh_op_bnl_6')
// (28, 20, 'sp4_h_l_41')

wire n166;
// (21, 17, 'neigh_op_tnr_0')
// (21, 18, 'neigh_op_rgt_0')
// (21, 19, 'local_g0_0')
// (21, 19, 'lutff_2/in_2')
// (21, 19, 'neigh_op_bnr_0')
// (22, 17, 'neigh_op_top_0')
// (22, 18, 'lutff_0/out')
// (22, 19, 'local_g0_0')
// (22, 19, 'lutff_2/in_2')
// (22, 19, 'neigh_op_bot_0')
// (23, 17, 'neigh_op_tnl_0')
// (23, 18, 'neigh_op_lft_0')
// (23, 19, 'neigh_op_bnl_0')

wire n167;
// (21, 17, 'neigh_op_tnr_2')
// (21, 18, 'neigh_op_rgt_2')
// (21, 19, 'local_g1_2')
// (21, 19, 'lutff_3/in_2')
// (21, 19, 'neigh_op_bnr_2')
// (22, 17, 'neigh_op_top_2')
// (22, 18, 'lutff_2/out')
// (22, 19, 'local_g1_2')
// (22, 19, 'lutff_3/in_2')
// (22, 19, 'neigh_op_bot_2')
// (23, 17, 'neigh_op_tnl_2')
// (23, 18, 'neigh_op_lft_2')
// (23, 19, 'neigh_op_bnl_2')

wire n168;
// (21, 17, 'neigh_op_tnr_5')
// (21, 18, 'neigh_op_rgt_5')
// (21, 19, 'local_g0_5')
// (21, 19, 'lutff_6/in_1')
// (21, 19, 'neigh_op_bnr_5')
// (22, 17, 'neigh_op_top_5')
// (22, 18, 'lutff_5/out')
// (22, 19, 'local_g1_5')
// (22, 19, 'lutff_6/in_2')
// (22, 19, 'neigh_op_bot_5')
// (23, 17, 'neigh_op_tnl_5')
// (23, 18, 'neigh_op_lft_5')
// (23, 19, 'neigh_op_bnl_5')

wire n169;
// (21, 17, 'neigh_op_tnr_7')
// (21, 18, 'neigh_op_rgt_7')
// (21, 19, 'local_g0_7')
// (21, 19, 'lutff_0/in_1')
// (21, 19, 'neigh_op_bnr_7')
// (22, 17, 'neigh_op_top_7')
// (22, 18, 'lutff_7/out')
// (22, 19, 'local_g0_7')
// (22, 19, 'lutff_0/in_1')
// (22, 19, 'neigh_op_bot_7')
// (23, 17, 'neigh_op_tnl_7')
// (23, 18, 'neigh_op_lft_7')
// (23, 19, 'neigh_op_bnl_7')

wire n170;
// (21, 19, 'lutff_7/cout')
// (21, 20, 'carry_in')
// (21, 20, 'carry_in_mux')

wire n171;
// (21, 20, 'local_g0_1')
// (21, 20, 'lutff_6/in_1')
// (21, 20, 'sp4_h_r_9')
// (22, 20, 'local_g0_4')
// (22, 20, 'lutff_6/in_2')
// (22, 20, 'sp4_h_r_20')
// (23, 19, 'neigh_op_tnr_6')
// (23, 20, 'neigh_op_rgt_6')
// (23, 20, 'sp4_h_r_33')
// (23, 21, 'neigh_op_bnr_6')
// (24, 19, 'neigh_op_top_6')
// (24, 20, 'lutff_6/out')
// (24, 20, 'sp4_h_r_44')
// (24, 21, 'neigh_op_bot_6')
// (25, 19, 'neigh_op_tnl_6')
// (25, 20, 'neigh_op_lft_6')
// (25, 20, 'sp4_h_l_44')
// (25, 21, 'neigh_op_bnl_6')

wire n172;
// (21, 20, 'local_g1_4')
// (21, 20, 'lutff_3/in_2')
// (21, 20, 'sp4_h_r_4')
// (22, 19, 'neigh_op_tnr_6')
// (22, 20, 'local_g3_6')
// (22, 20, 'lutff_3/in_2')
// (22, 20, 'neigh_op_rgt_6')
// (22, 20, 'sp4_h_r_17')
// (22, 21, 'neigh_op_bnr_6')
// (23, 19, 'neigh_op_top_6')
// (23, 20, 'lutff_6/out')
// (23, 20, 'sp4_h_r_28')
// (23, 21, 'neigh_op_bot_6')
// (24, 19, 'neigh_op_tnl_6')
// (24, 20, 'neigh_op_lft_6')
// (24, 20, 'sp4_h_r_41')
// (24, 21, 'neigh_op_bnl_6')
// (25, 20, 'sp4_h_l_41')

wire n173;
// (21, 20, 'local_g2_3')
// (21, 20, 'lutff_2/in_1')
// (21, 20, 'neigh_op_tnr_3')
// (21, 21, 'neigh_op_rgt_3')
// (21, 22, 'neigh_op_bnr_3')
// (22, 20, 'local_g1_3')
// (22, 20, 'lutff_2/in_2')
// (22, 20, 'neigh_op_top_3')
// (22, 21, 'lutff_3/out')
// (22, 22, 'neigh_op_bot_3')
// (23, 20, 'neigh_op_tnl_3')
// (23, 21, 'neigh_op_lft_3')
// (23, 22, 'neigh_op_bnl_3')

wire n174;
// (21, 20, 'local_g2_6')
// (21, 20, 'lutff_5/in_1')
// (21, 20, 'neigh_op_tnr_6')
// (21, 21, 'neigh_op_rgt_6')
// (21, 22, 'neigh_op_bnr_6')
// (22, 20, 'local_g0_6')
// (22, 20, 'lutff_5/in_1')
// (22, 20, 'neigh_op_top_6')
// (22, 21, 'lutff_6/out')
// (22, 22, 'neigh_op_bot_6')
// (23, 20, 'neigh_op_tnl_6')
// (23, 21, 'neigh_op_lft_6')
// (23, 22, 'neigh_op_bnl_6')

wire n175;
// (21, 20, 'local_g3_5')
// (21, 20, 'lutff_0/in_2')
// (21, 20, 'neigh_op_tnr_5')
// (21, 21, 'neigh_op_rgt_5')
// (21, 22, 'neigh_op_bnr_5')
// (22, 20, 'local_g0_5')
// (22, 20, 'lutff_0/in_1')
// (22, 20, 'neigh_op_top_5')
// (22, 21, 'lutff_5/out')
// (22, 22, 'neigh_op_bot_5')
// (23, 20, 'neigh_op_tnl_5')
// (23, 21, 'neigh_op_lft_5')
// (23, 22, 'neigh_op_bnl_5')

wire n176;
// (21, 20, 'lutff_7/cout')
// (21, 21, 'carry_in')
// (21, 21, 'carry_in_mux')
// (21, 21, 'lutff_0/in_3')

wire n177;
// (21, 20, 'neigh_op_tnr_0')
// (21, 21, 'neigh_op_rgt_0')
// (21, 22, 'neigh_op_bnr_0')
// (22, 20, 'neigh_op_top_0')
// (22, 21, 'local_g0_0')
// (22, 21, 'lutff_0/out')
// (22, 21, 'lutff_4/in_0')
// (22, 22, 'neigh_op_bot_0')
// (23, 20, 'neigh_op_tnl_0')
// (23, 21, 'neigh_op_lft_0')
// (23, 22, 'neigh_op_bnl_0')

wire n178;
// (21, 21, 'neigh_op_tnr_6')
// (21, 22, 'neigh_op_rgt_6')
// (21, 23, 'neigh_op_bnr_6')
// (22, 21, 'neigh_op_top_6')
// (22, 22, 'lutff_6/out')
// (22, 23, 'neigh_op_bot_6')
// (23, 21, 'local_g2_6')
// (23, 21, 'lutff_0/in_0')
// (23, 21, 'neigh_op_tnl_6')
// (23, 22, 'neigh_op_lft_6')
// (23, 23, 'neigh_op_bnl_6')

wire n179;
// (21, 21, 'sp4_h_r_1')
// (22, 21, 'local_g1_4')
// (22, 21, 'lutff_4/in_3')
// (22, 21, 'sp4_h_r_12')
// (23, 20, 'neigh_op_tnr_2')
// (23, 21, 'neigh_op_rgt_2')
// (23, 21, 'sp4_h_r_25')
// (23, 22, 'neigh_op_bnr_2')
// (24, 20, 'neigh_op_top_2')
// (24, 21, 'lutff_2/out')
// (24, 21, 'sp4_h_r_36')
// (24, 22, 'neigh_op_bot_2')
// (25, 20, 'neigh_op_tnl_2')
// (25, 21, 'neigh_op_lft_2')
// (25, 21, 'sp4_h_l_36')
// (25, 22, 'neigh_op_bnl_2')

wire io_33_23_1;
// (22, 11, 'sp12_v_t_23')
// (22, 12, 'sp12_v_b_23')
// (22, 13, 'sp12_v_b_20')
// (22, 14, 'sp12_v_b_19')
// (22, 15, 'sp12_v_b_16')
// (22, 16, 'sp12_v_b_15')
// (22, 17, 'sp12_v_b_12')
// (22, 18, 'sp12_v_b_11')
// (22, 19, 'sp12_v_b_8')
// (22, 20, 'sp12_v_b_7')
// (22, 21, 'local_g2_4')
// (22, 21, 'lutff_4/in_2')
// (22, 21, 'lutff_6/in_2')
// (22, 21, 'sp12_v_b_4')
// (22, 22, 'sp12_v_b_3')
// (22, 23, 'sp12_h_r_0')
// (22, 23, 'sp12_v_b_0')
// (23, 23, 'sp12_h_r_3')
// (24, 23, 'sp12_h_r_4')
// (25, 23, 'sp12_h_r_7')
// (26, 23, 'sp12_h_r_8')
// (27, 23, 'sp12_h_r_11')
// (28, 23, 'sp12_h_r_12')
// (29, 23, 'sp12_h_r_15')
// (30, 23, 'sp12_h_r_16')
// (31, 23, 'sp12_h_r_19')
// (32, 22, 'neigh_op_tnr_2')
// (32, 22, 'neigh_op_tnr_6')
// (32, 23, 'neigh_op_rgt_2')
// (32, 23, 'neigh_op_rgt_6')
// (32, 23, 'sp12_h_r_20')
// (32, 24, 'neigh_op_bnr_2')
// (32, 24, 'neigh_op_bnr_6')
// (33, 23, 'io_1/D_IN_0')
// (33, 23, 'io_1/PAD')
// (33, 23, 'span12_horz_20')

wire n181;
// (22, 19, 'lutff_7/cout')
// (22, 20, 'carry_in')
// (22, 20, 'carry_in_mux')

wire n182;
// (22, 20, 'lutff_7/cout')
// (22, 21, 'carry_in')
// (22, 21, 'carry_in_mux')
// (22, 21, 'lutff_0/in_3')

wire n183;
// (22, 20, 'neigh_op_tnr_0')
// (22, 21, 'neigh_op_rgt_0')
// (22, 22, 'neigh_op_bnr_0')
// (23, 20, 'neigh_op_top_0')
// (23, 21, 'local_g0_0')
// (23, 21, 'lutff_0/out')
// (23, 21, 'lutff_1/in_1')
// (23, 22, 'neigh_op_bot_0')
// (24, 20, 'neigh_op_tnl_0')
// (24, 21, 'neigh_op_lft_0')
// (24, 22, 'neigh_op_bnl_0')

wire n184;
// (22, 20, 'neigh_op_tnr_1')
// (22, 21, 'local_g2_1')
// (22, 21, 'lutff_4/in_1')
// (22, 21, 'neigh_op_rgt_1')
// (22, 22, 'neigh_op_bnr_1')
// (23, 20, 'neigh_op_top_1')
// (23, 21, 'lutff_1/out')
// (23, 22, 'neigh_op_bot_1')
// (24, 20, 'neigh_op_tnl_1')
// (24, 21, 'neigh_op_lft_1')
// (24, 22, 'neigh_op_bnl_1')

wire n185;
// (22, 20, 'neigh_op_tnr_6')
// (22, 21, 'neigh_op_rgt_6')
// (22, 22, 'neigh_op_bnr_6')
// (23, 20, 'neigh_op_top_6')
// (23, 21, 'local_g0_6')
// (23, 21, 'lutff_1/in_3')
// (23, 21, 'lutff_6/out')
// (23, 22, 'neigh_op_bot_6')
// (24, 20, 'neigh_op_tnl_6')
// (24, 21, 'neigh_op_lft_6')
// (24, 22, 'neigh_op_bnl_6')

wire io_33_20_1;
// (22, 20, 'sp12_h_r_0')
// (23, 20, 'sp12_h_r_3')
// (24, 19, 'sp4_r_v_b_37')
// (24, 20, 'local_g0_4')
// (24, 20, 'lutff_6/in_2')
// (24, 20, 'sp12_h_r_4')
// (24, 20, 'sp4_r_v_b_24')
// (24, 21, 'local_g2_5')
// (24, 21, 'lutff_2/in_3')
// (24, 21, 'sp4_r_v_b_13')
// (24, 22, 'sp4_r_v_b_0')
// (25, 18, 'sp4_v_t_37')
// (25, 19, 'sp4_v_b_37')
// (25, 20, 'sp12_h_r_7')
// (25, 20, 'sp4_v_b_24')
// (25, 21, 'sp4_v_b_13')
// (25, 22, 'sp4_h_r_0')
// (25, 22, 'sp4_v_b_0')
// (26, 20, 'sp12_h_r_8')
// (26, 22, 'sp4_h_r_13')
// (27, 20, 'sp12_h_r_11')
// (27, 22, 'sp4_h_r_24')
// (28, 20, 'sp12_h_r_12')
// (28, 22, 'sp4_h_r_37')
// (29, 20, 'sp12_h_r_15')
// (29, 22, 'sp4_h_l_37')
// (29, 22, 'sp4_h_r_0')
// (30, 20, 'sp12_h_r_16')
// (30, 22, 'sp4_h_r_13')
// (31, 20, 'sp12_h_r_19')
// (31, 22, 'sp4_h_r_24')
// (32, 19, 'neigh_op_tnr_2')
// (32, 19, 'neigh_op_tnr_6')
// (32, 20, 'neigh_op_rgt_2')
// (32, 20, 'neigh_op_rgt_6')
// (32, 20, 'sp12_h_r_20')
// (32, 21, 'neigh_op_bnr_2')
// (32, 21, 'neigh_op_bnr_6')
// (32, 22, 'sp4_h_r_37')
// (33, 18, 'span4_vert_t_14')
// (33, 19, 'span4_vert_b_14')
// (33, 20, 'io_1/D_IN_0')
// (33, 20, 'io_1/PAD')
// (33, 20, 'span12_horz_20')
// (33, 20, 'span4_vert_b_10')
// (33, 21, 'span4_vert_b_6')
// (33, 22, 'span4_horz_37')
// (33, 22, 'span4_vert_b_2')

wire io_33_21_1;
// (22, 21, 'sp12_h_r_0')
// (23, 18, 'sp4_r_v_b_38')
// (23, 19, 'sp4_r_v_b_27')
// (23, 20, 'local_g2_6')
// (23, 20, 'lutff_2/in_2')
// (23, 20, 'lutff_4/in_0')
// (23, 20, 'sp4_r_v_b_14')
// (23, 21, 'sp12_h_r_3')
// (23, 21, 'sp4_r_v_b_3')
// (24, 17, 'sp4_v_t_38')
// (24, 18, 'sp4_r_v_b_47')
// (24, 18, 'sp4_v_b_38')
// (24, 19, 'sp4_r_v_b_34')
// (24, 19, 'sp4_v_b_27')
// (24, 20, 'local_g3_7')
// (24, 20, 'lutff_1/in_1')
// (24, 20, 'sp4_r_v_b_23')
// (24, 20, 'sp4_v_b_14')
// (24, 21, 'local_g1_4')
// (24, 21, 'lutff_4/in_1')
// (24, 21, 'sp12_h_r_4')
// (24, 21, 'sp4_h_r_3')
// (24, 21, 'sp4_r_v_b_10')
// (24, 21, 'sp4_v_b_3')
// (25, 17, 'sp4_v_t_47')
// (25, 18, 'sp4_r_v_b_41')
// (25, 18, 'sp4_v_b_47')
// (25, 19, 'sp4_r_v_b_28')
// (25, 19, 'sp4_v_b_34')
// (25, 20, 'sp4_r_v_b_17')
// (25, 20, 'sp4_v_b_23')
// (25, 21, 'sp12_h_r_7')
// (25, 21, 'sp4_h_r_14')
// (25, 21, 'sp4_h_r_5')
// (25, 21, 'sp4_r_v_b_4')
// (25, 21, 'sp4_v_b_10')
// (26, 17, 'sp4_v_t_41')
// (26, 18, 'sp4_v_b_41')
// (26, 19, 'sp4_v_b_28')
// (26, 20, 'local_g1_1')
// (26, 20, 'lutff_6/in_0')
// (26, 20, 'sp4_v_b_17')
// (26, 21, 'local_g1_0')
// (26, 21, 'lutff_2/in_1')
// (26, 21, 'sp12_h_r_0')
// (26, 21, 'sp12_h_r_8')
// (26, 21, 'sp4_h_r_16')
// (26, 21, 'sp4_h_r_27')
// (26, 21, 'sp4_h_r_4')
// (26, 21, 'sp4_v_b_4')
// (27, 21, 'sp12_h_r_11')
// (27, 21, 'sp12_h_r_3')
// (27, 21, 'sp4_h_r_17')
// (27, 21, 'sp4_h_r_29')
// (27, 21, 'sp4_h_r_38')
// (28, 21, 'sp12_h_r_12')
// (28, 21, 'sp12_h_r_4')
// (28, 21, 'sp4_h_l_38')
// (28, 21, 'sp4_h_r_0')
// (28, 21, 'sp4_h_r_28')
// (28, 21, 'sp4_h_r_40')
// (29, 21, 'sp12_h_r_15')
// (29, 21, 'sp12_h_r_7')
// (29, 21, 'sp4_h_l_40')
// (29, 21, 'sp4_h_r_13')
// (29, 21, 'sp4_h_r_41')
// (29, 21, 'sp4_h_r_9')
// (30, 21, 'sp12_h_r_16')
// (30, 21, 'sp12_h_r_8')
// (30, 21, 'sp4_h_l_41')
// (30, 21, 'sp4_h_r_20')
// (30, 21, 'sp4_h_r_24')
// (30, 21, 'sp4_h_r_4')
// (31, 21, 'sp12_h_r_11')
// (31, 21, 'sp12_h_r_19')
// (31, 21, 'sp4_h_r_17')
// (31, 21, 'sp4_h_r_33')
// (31, 21, 'sp4_h_r_37')
// (32, 20, 'neigh_op_tnr_2')
// (32, 20, 'neigh_op_tnr_6')
// (32, 21, 'neigh_op_rgt_2')
// (32, 21, 'neigh_op_rgt_6')
// (32, 21, 'sp12_h_r_12')
// (32, 21, 'sp12_h_r_20')
// (32, 21, 'sp4_h_l_37')
// (32, 21, 'sp4_h_r_28')
// (32, 21, 'sp4_h_r_4')
// (32, 21, 'sp4_h_r_44')
// (32, 22, 'neigh_op_bnr_2')
// (32, 22, 'neigh_op_bnr_6')
// (33, 21, 'io_1/D_IN_0')
// (33, 21, 'io_1/PAD')
// (33, 21, 'span12_horz_12')
// (33, 21, 'span12_horz_20')
// (33, 21, 'span4_horz_28')
// (33, 21, 'span4_horz_4')
// (33, 21, 'span4_horz_44')

wire io_33_28_0;
// (23, 17, 'sp4_r_v_b_45')
// (23, 18, 'sp4_r_v_b_32')
// (23, 19, 'sp4_r_v_b_21')
// (23, 20, 'local_g2_0')
// (23, 20, 'lutff_2/in_0')
// (23, 20, 'lutff_4/in_2')
// (23, 20, 'lutff_6/in_0')
// (23, 20, 'sp4_r_v_b_8')
// (24, 16, 'sp12_v_t_23')
// (24, 16, 'sp4_v_t_45')
// (24, 17, 'sp12_v_b_23')
// (24, 17, 'sp4_v_b_45')
// (24, 18, 'sp12_v_b_20')
// (24, 18, 'sp4_v_b_32')
// (24, 19, 'sp12_v_b_19')
// (24, 19, 'sp4_v_b_21')
// (24, 20, 'local_g3_0')
// (24, 20, 'lutff_1/in_0')
// (24, 20, 'sp12_v_b_16')
// (24, 20, 'sp4_v_b_8')
// (24, 21, 'local_g3_7')
// (24, 21, 'lutff_4/in_2')
// (24, 21, 'sp12_v_b_15')
// (24, 22, 'sp12_v_b_12')
// (24, 23, 'sp12_v_b_11')
// (24, 24, 'sp12_v_b_8')
// (24, 25, 'sp12_v_b_7')
// (24, 26, 'sp12_v_b_4')
// (24, 27, 'sp12_v_b_3')
// (24, 28, 'sp12_h_r_0')
// (24, 28, 'sp12_v_b_0')
// (25, 28, 'sp12_h_r_3')
// (26, 21, 'local_g1_1')
// (26, 21, 'lutff_2/in_2')
// (26, 21, 'sp4_h_r_9')
// (26, 28, 'sp12_h_r_4')
// (27, 21, 'sp4_h_r_20')
// (27, 28, 'sp12_h_r_7')
// (28, 21, 'sp4_h_r_33')
// (28, 28, 'sp12_h_r_8')
// (29, 21, 'sp4_h_r_44')
// (29, 28, 'sp12_h_r_11')
// (30, 21, 'sp4_h_l_44')
// (30, 21, 'sp4_h_r_1')
// (30, 28, 'sp12_h_r_12')
// (31, 21, 'sp4_h_r_12')
// (31, 28, 'sp12_h_r_15')
// (32, 21, 'sp4_h_r_25')
// (32, 27, 'neigh_op_tnr_0')
// (32, 27, 'neigh_op_tnr_4')
// (32, 28, 'neigh_op_rgt_0')
// (32, 28, 'neigh_op_rgt_4')
// (32, 28, 'sp12_h_r_16')
// (32, 29, 'neigh_op_bnr_0')
// (32, 29, 'neigh_op_bnr_4')
// (33, 21, 'span4_horz_25')
// (33, 21, 'span4_vert_t_12')
// (33, 22, 'span4_vert_b_12')
// (33, 23, 'span4_vert_b_8')
// (33, 24, 'span4_vert_b_4')
// (33, 25, 'span4_vert_b_0')
// (33, 25, 'span4_vert_t_12')
// (33, 26, 'span4_vert_b_12')
// (33, 27, 'span4_vert_b_8')
// (33, 28, 'io_0/D_IN_0')
// (33, 28, 'io_0/PAD')
// (33, 28, 'span12_horz_16')
// (33, 28, 'span4_vert_b_4')
// (33, 29, 'span4_vert_b_0')

wire n189;
// (23, 20, 'neigh_op_tnr_4')
// (23, 20, 'sp4_r_v_b_37')
// (23, 21, 'neigh_op_rgt_4')
// (23, 21, 'sp4_r_v_b_24')
// (23, 22, 'neigh_op_bnr_4')
// (23, 22, 'sp4_r_v_b_13')
// (23, 23, 'sp4_r_v_b_0')
// (24, 17, 'sp4_r_v_b_42')
// (24, 18, 'sp4_r_v_b_31')
// (24, 18, 'sp4_r_v_b_44')
// (24, 19, 'sp4_r_v_b_18')
// (24, 19, 'sp4_r_v_b_33')
// (24, 19, 'sp4_v_t_37')
// (24, 20, 'neigh_op_top_4')
// (24, 20, 'sp4_r_v_b_20')
// (24, 20, 'sp4_r_v_b_7')
// (24, 20, 'sp4_v_b_37')
// (24, 21, 'lutff_4/out')
// (24, 21, 'sp4_r_v_b_41')
// (24, 21, 'sp4_r_v_b_9')
// (24, 21, 'sp4_v_b_24')
// (24, 22, 'local_g0_4')
// (24, 22, 'lutff_5/in_1')
// (24, 22, 'neigh_op_bot_4')
// (24, 22, 'sp4_r_v_b_28')
// (24, 22, 'sp4_v_b_13')
// (24, 23, 'sp4_h_r_6')
// (24, 23, 'sp4_r_v_b_17')
// (24, 23, 'sp4_v_b_0')
// (24, 24, 'sp4_r_v_b_4')
// (24, 25, 'sp4_r_v_b_42')
// (24, 26, 'sp4_r_v_b_31')
// (24, 27, 'sp4_r_v_b_18')
// (24, 28, 'sp4_r_v_b_7')
// (25, 16, 'sp4_v_t_42')
// (25, 17, 'local_g0_2')
// (25, 17, 'ram/RCLKE')
// (25, 17, 'sp4_h_r_2')
// (25, 17, 'sp4_v_b_42')
// (25, 17, 'sp4_v_t_44')
// (25, 18, 'sp4_v_b_31')
// (25, 18, 'sp4_v_b_44')
// (25, 19, 'local_g0_2')
// (25, 19, 'ram/RCLKE')
// (25, 19, 'sp4_v_b_18')
// (25, 19, 'sp4_v_b_33')
// (25, 20, 'neigh_op_tnl_4')
// (25, 20, 'sp4_v_b_20')
// (25, 20, 'sp4_v_b_7')
// (25, 20, 'sp4_v_t_41')
// (25, 21, 'neigh_op_lft_4')
// (25, 21, 'sp4_v_b_41')
// (25, 21, 'sp4_v_b_9')
// (25, 22, 'neigh_op_bnl_4')
// (25, 22, 'sp4_v_b_28')
// (25, 23, 'local_g1_3')
// (25, 23, 'ram/RCLKE')
// (25, 23, 'sp4_h_r_19')
// (25, 23, 'sp4_v_b_17')
// (25, 24, 'sp4_v_b_4')
// (25, 24, 'sp4_v_t_42')
// (25, 25, 'sp4_v_b_42')
// (25, 26, 'sp4_v_b_31')
// (25, 27, 'local_g0_2')
// (25, 27, 'ram/RCLKE')
// (25, 27, 'sp4_v_b_18')
// (25, 28, 'sp4_v_b_7')
// (26, 17, 'sp4_h_r_15')
// (26, 23, 'sp4_h_r_30')
// (27, 17, 'sp4_h_r_26')
// (27, 23, 'sp4_h_r_43')
// (28, 17, 'sp4_h_r_39')
// (28, 23, 'sp4_h_l_43')
// (29, 17, 'sp4_h_l_39')

wire n190;
// (23, 21, 'sp4_h_r_1')
// (24, 21, 'local_g0_4')
// (24, 21, 'lutff_2/in_0')
// (24, 21, 'sp4_h_r_12')
// (25, 20, 'neigh_op_tnr_2')
// (25, 21, 'neigh_op_rgt_2')
// (25, 21, 'sp4_h_r_25')
// (25, 22, 'neigh_op_bnr_2')
// (26, 20, 'neigh_op_top_2')
// (26, 21, 'lutff_2/out')
// (26, 21, 'sp4_h_r_36')
// (26, 22, 'neigh_op_bot_2')
// (27, 20, 'neigh_op_tnl_2')
// (27, 21, 'neigh_op_lft_2')
// (27, 21, 'sp4_h_l_36')
// (27, 22, 'neigh_op_bnl_2')

wire n191;
// (23, 25, 'neigh_op_tnr_0')
// (23, 26, 'neigh_op_rgt_0')
// (23, 27, 'neigh_op_bnr_0')
// (24, 25, 'local_g1_0')
// (24, 25, 'lutff_5/in_2')
// (24, 25, 'neigh_op_top_0')
// (24, 26, 'lutff_0/out')
// (24, 27, 'neigh_op_bot_0')
// (25, 25, 'neigh_op_tnl_0')
// (25, 26, 'neigh_op_lft_0')
// (25, 27, 'neigh_op_bnl_0')

wire n192;
// (23, 25, 'neigh_op_tnr_1')
// (23, 26, 'neigh_op_rgt_1')
// (23, 27, 'neigh_op_bnr_1')
// (24, 25, 'local_g1_1')
// (24, 25, 'lutff_7/in_3')
// (24, 25, 'neigh_op_top_1')
// (24, 26, 'lutff_1/out')
// (24, 27, 'neigh_op_bot_1')
// (25, 25, 'neigh_op_tnl_1')
// (25, 26, 'neigh_op_lft_1')
// (25, 27, 'neigh_op_bnl_1')

wire n193;
// (24, 14, 'neigh_op_tnr_4')
// (24, 14, 'sp4_r_v_b_37')
// (24, 15, 'neigh_op_rgt_4')
// (24, 15, 'sp4_r_v_b_24')
// (24, 16, 'neigh_op_bnr_4')
// (24, 16, 'sp4_r_v_b_13')
// (24, 17, 'local_g1_0')
// (24, 17, 'lutff_5/in_2')
// (24, 17, 'sp4_r_v_b_0')
// (25, 13, 'sp4_v_t_37')
// (25, 14, 'neigh_op_top_4')
// (25, 14, 'sp4_v_b_37')
// (25, 15, 'ram/RDATA_11')
// (25, 15, 'sp4_v_b_24')
// (25, 16, 'neigh_op_bot_4')
// (25, 16, 'sp4_v_b_13')
// (25, 17, 'sp4_v_b_0')
// (26, 14, 'neigh_op_tnl_4')
// (26, 15, 'neigh_op_lft_4')
// (26, 16, 'neigh_op_bnl_4')

wire n194;
// (24, 15, 'neigh_op_tnr_4')
// (24, 16, 'neigh_op_rgt_4')
// (24, 17, 'local_g0_4')
// (24, 17, 'lutff_7/in_3')
// (24, 17, 'neigh_op_bnr_4')
// (25, 15, 'neigh_op_top_4')
// (25, 16, 'ram/RDATA_3')
// (25, 17, 'neigh_op_bot_4')
// (26, 15, 'neigh_op_tnl_4')
// (26, 16, 'neigh_op_lft_4')
// (26, 17, 'neigh_op_bnl_4')

wire n195;
// (24, 16, 'neigh_op_tnr_4')
// (24, 17, 'local_g2_4')
// (24, 17, 'lutff_5/in_3')
// (24, 17, 'neigh_op_rgt_4')
// (24, 18, 'neigh_op_bnr_4')
// (25, 16, 'neigh_op_top_4')
// (25, 17, 'ram/RDATA_11')
// (25, 18, 'neigh_op_bot_4')
// (26, 16, 'neigh_op_tnl_4')
// (26, 17, 'neigh_op_lft_4')
// (26, 18, 'neigh_op_bnl_4')

wire n196;
// (24, 17, 'local_g3_4')
// (24, 17, 'lutff_7/in_0')
// (24, 17, 'neigh_op_tnr_4')
// (24, 18, 'neigh_op_rgt_4')
// (24, 19, 'neigh_op_bnr_4')
// (25, 17, 'neigh_op_top_4')
// (25, 18, 'ram/RDATA_3')
// (25, 19, 'neigh_op_bot_4')
// (26, 17, 'neigh_op_tnl_4')
// (26, 18, 'neigh_op_lft_4')
// (26, 19, 'neigh_op_bnl_4')

wire n197;
// (24, 20, 'neigh_op_tnr_4')
// (24, 21, 'local_g3_4')
// (24, 21, 'lutff_7/in_2')
// (24, 21, 'neigh_op_rgt_4')
// (24, 22, 'neigh_op_bnr_4')
// (25, 20, 'neigh_op_top_4')
// (25, 21, 'ram/RDATA_11')
// (25, 22, 'neigh_op_bot_4')
// (26, 20, 'neigh_op_tnl_4')
// (26, 21, 'neigh_op_lft_4')
// (26, 22, 'neigh_op_bnl_4')

wire n198;
// (24, 20, 'sp4_r_v_b_45')
// (24, 21, 'local_g0_3')
// (24, 21, 'lutff_7/in_0')
// (24, 21, 'sp4_r_v_b_32')
// (24, 22, 'neigh_op_tnr_4')
// (24, 22, 'sp4_r_v_b_21')
// (24, 23, 'neigh_op_rgt_4')
// (24, 23, 'sp4_r_v_b_8')
// (24, 24, 'neigh_op_bnr_4')
// (25, 19, 'sp4_v_t_45')
// (25, 20, 'sp4_v_b_45')
// (25, 21, 'sp4_v_b_32')
// (25, 22, 'neigh_op_top_4')
// (25, 22, 'sp4_v_b_21')
// (25, 23, 'ram/RDATA_11')
// (25, 23, 'sp4_v_b_8')
// (25, 24, 'neigh_op_bot_4')
// (26, 22, 'neigh_op_tnl_4')
// (26, 23, 'neigh_op_lft_4')
// (26, 24, 'neigh_op_bnl_4')

wire io_33_21_0;
// (24, 21, 'local_g0_0')
// (24, 21, 'local_g1_0')
// (24, 21, 'lutff_2/in_2')
// (24, 21, 'lutff_3/in_0')
// (24, 21, 'sp12_h_r_0')
// (25, 21, 'sp12_h_r_3')
// (26, 21, 'sp12_h_r_4')
// (27, 21, 'sp12_h_r_7')
// (28, 21, 'sp12_h_r_8')
// (29, 21, 'sp12_h_r_11')
// (30, 21, 'sp12_h_r_12')
// (31, 21, 'sp12_h_r_15')
// (32, 20, 'neigh_op_tnr_0')
// (32, 20, 'neigh_op_tnr_4')
// (32, 21, 'neigh_op_rgt_0')
// (32, 21, 'neigh_op_rgt_4')
// (32, 21, 'sp12_h_r_16')
// (32, 22, 'neigh_op_bnr_0')
// (32, 22, 'neigh_op_bnr_4')
// (33, 21, 'io_0/D_IN_0')
// (33, 21, 'io_0/PAD')
// (33, 21, 'span12_horz_16')

wire n200;
// (24, 21, 'neigh_op_tnr_4')
// (24, 22, 'local_g2_4')
// (24, 22, 'lutff_7/in_1')
// (24, 22, 'neigh_op_rgt_4')
// (24, 23, 'neigh_op_bnr_4')
// (25, 21, 'neigh_op_top_4')
// (25, 22, 'ram/RDATA_3')
// (25, 23, 'neigh_op_bot_4')
// (26, 21, 'neigh_op_tnl_4')
// (26, 22, 'neigh_op_lft_4')
// (26, 23, 'neigh_op_bnl_4')

wire n201;
// (24, 21, 'sp4_r_v_b_45')
// (24, 22, 'local_g0_3')
// (24, 22, 'lutff_7/in_2')
// (24, 22, 'sp4_r_v_b_32')
// (24, 23, 'neigh_op_tnr_4')
// (24, 23, 'sp4_r_v_b_21')
// (24, 24, 'neigh_op_rgt_4')
// (24, 24, 'sp4_r_v_b_8')
// (24, 25, 'neigh_op_bnr_4')
// (25, 20, 'sp4_v_t_45')
// (25, 21, 'sp4_v_b_45')
// (25, 22, 'sp4_v_b_32')
// (25, 23, 'neigh_op_top_4')
// (25, 23, 'sp4_v_b_21')
// (25, 24, 'ram/RDATA_3')
// (25, 24, 'sp4_v_b_8')
// (25, 25, 'neigh_op_bot_4')
// (26, 23, 'neigh_op_tnl_4')
// (26, 24, 'neigh_op_lft_4')
// (26, 25, 'neigh_op_bnl_4')

wire n202;
// (24, 23, 'sp4_r_v_b_41')
// (24, 24, 'sp4_r_v_b_28')
// (24, 25, 'sp4_r_v_b_17')
// (24, 26, 'local_g1_4')
// (24, 26, 'lutff_0/in_3')
// (24, 26, 'sp4_r_v_b_4')
// (24, 27, 'sp4_r_v_b_45')
// (24, 28, 'sp4_r_v_b_32')
// (24, 29, 'neigh_op_tnr_4')
// (24, 29, 'sp4_r_v_b_21')
// (24, 30, 'neigh_op_rgt_4')
// (24, 30, 'sp4_r_v_b_8')
// (24, 31, 'neigh_op_bnr_4')
// (25, 22, 'sp4_v_t_41')
// (25, 23, 'sp4_v_b_41')
// (25, 24, 'sp4_v_b_28')
// (25, 25, 'sp4_v_b_17')
// (25, 26, 'sp4_v_b_4')
// (25, 26, 'sp4_v_t_45')
// (25, 27, 'sp4_v_b_45')
// (25, 28, 'sp4_v_b_32')
// (25, 29, 'neigh_op_top_4')
// (25, 29, 'sp4_v_b_21')
// (25, 30, 'ram/RDATA_3')
// (25, 30, 'sp4_v_b_8')
// (25, 31, 'neigh_op_bot_4')
// (26, 29, 'neigh_op_tnl_4')
// (26, 30, 'neigh_op_lft_4')
// (26, 31, 'neigh_op_bnl_4')

wire n203;
// (24, 24, 'neigh_op_tnr_4')
// (24, 25, 'local_g3_4')
// (24, 25, 'lutff_7/in_0')
// (24, 25, 'neigh_op_rgt_4')
// (24, 26, 'neigh_op_bnr_4')
// (25, 24, 'neigh_op_top_4')
// (25, 25, 'ram/RDATA_11')
// (25, 26, 'neigh_op_bot_4')
// (26, 24, 'neigh_op_tnl_4')
// (26, 25, 'neigh_op_lft_4')
// (26, 26, 'neigh_op_bnl_4')

wire n204;
// (24, 25, 'local_g2_4')
// (24, 25, 'lutff_5/in_3')
// (24, 25, 'neigh_op_tnr_4')
// (24, 26, 'neigh_op_rgt_4')
// (24, 27, 'neigh_op_bnr_4')
// (25, 25, 'neigh_op_top_4')
// (25, 26, 'ram/RDATA_3')
// (25, 27, 'neigh_op_bot_4')
// (26, 25, 'neigh_op_tnl_4')
// (26, 26, 'neigh_op_lft_4')
// (26, 27, 'neigh_op_bnl_4')

wire n205;
// (24, 25, 'sp4_r_v_b_45')
// (24, 26, 'local_g2_0')
// (24, 26, 'lutff_0/in_0')
// (24, 26, 'sp4_r_v_b_32')
// (24, 27, 'neigh_op_tnr_4')
// (24, 27, 'sp4_r_v_b_21')
// (24, 28, 'neigh_op_rgt_4')
// (24, 28, 'sp4_r_v_b_8')
// (24, 29, 'neigh_op_bnr_4')
// (25, 24, 'sp4_v_t_45')
// (25, 25, 'sp4_v_b_45')
// (25, 26, 'sp4_v_b_32')
// (25, 27, 'neigh_op_top_4')
// (25, 27, 'sp4_v_b_21')
// (25, 28, 'ram/RDATA_3')
// (25, 28, 'sp4_v_b_8')
// (25, 29, 'neigh_op_bot_4')
// (26, 27, 'neigh_op_tnl_4')
// (26, 28, 'neigh_op_lft_4')
// (26, 29, 'neigh_op_bnl_4')

wire n206;
// (24, 26, 'local_g3_4')
// (24, 26, 'lutff_1/in_0')
// (24, 26, 'neigh_op_tnr_4')
// (24, 27, 'neigh_op_rgt_4')
// (24, 28, 'neigh_op_bnr_4')
// (25, 26, 'neigh_op_top_4')
// (25, 27, 'ram/RDATA_11')
// (25, 28, 'neigh_op_bot_4')
// (26, 26, 'neigh_op_tnl_4')
// (26, 27, 'neigh_op_lft_4')
// (26, 28, 'neigh_op_bnl_4')

wire n207;
// (24, 26, 'local_g3_5')
// (24, 26, 'lutff_1/in_3')
// (24, 26, 'sp4_r_v_b_45')
// (24, 27, 'sp4_r_v_b_32')
// (24, 28, 'neigh_op_tnr_4')
// (24, 28, 'sp4_r_v_b_21')
// (24, 29, 'neigh_op_rgt_4')
// (24, 29, 'sp4_r_v_b_8')
// (24, 30, 'neigh_op_bnr_4')
// (25, 25, 'sp4_v_t_45')
// (25, 26, 'sp4_v_b_45')
// (25, 27, 'sp4_v_b_32')
// (25, 28, 'neigh_op_top_4')
// (25, 28, 'sp4_v_b_21')
// (25, 29, 'ram/RDATA_11')
// (25, 29, 'sp4_v_b_8')
// (25, 30, 'neigh_op_bot_4')
// (26, 28, 'neigh_op_tnl_4')
// (26, 29, 'neigh_op_lft_4')
// (26, 30, 'neigh_op_bnl_4')

wire n208;
// (25, 18, 'neigh_op_tnr_7')
// (25, 19, 'local_g2_7')
// (25, 19, 'neigh_op_rgt_7')
// (25, 19, 'ram/RADDR_6')
// (25, 20, 'neigh_op_bnr_7')
// (26, 18, 'neigh_op_top_7')
// (26, 19, 'lutff_7/out')
// (26, 20, 'neigh_op_bot_7')
// (27, 18, 'neigh_op_tnl_7')
// (27, 19, 'neigh_op_lft_7')
// (27, 20, 'neigh_op_bnl_7')

wire io_31_0_1;
// (29, 0, 'logic_op_tnr_6')
// (29, 1, 'neigh_op_rgt_6')
// (29, 2, 'neigh_op_bnr_6')
// (30, 0, 'logic_op_top_6')
// (30, 1, 'lutff_6/out')
// (30, 2, 'neigh_op_bot_6')
// (31, 0, 'io_1/D_OUT_0')
// (31, 0, 'io_1/PAD')
// (31, 0, 'local_g1_6')
// (31, 0, 'logic_op_tnl_6')
// (31, 1, 'neigh_op_lft_6')
// (31, 2, 'neigh_op_bnl_6')

wire open_0;
wire open_1;
wire open_2;
wire open_3;
wire open_4;
wire open_5;
wire open_6;
wire open_7;
wire open_8;
wire open_9;
wire open_10;
wire open_11;
wire open_12;
wire open_13;
wire open_14;
wire open_15;
wire open_16;
wire open_17;
wire open_18;
wire open_19;
wire open_20;
wire open_21;
wire open_22;
wire open_23;
wire open_24;
wire open_25;
wire open_26;
wire open_27;
wire open_28;
wire open_29;
wire open_30;
wire open_31;
wire open_32;
wire open_33;
wire open_34;
wire open_35;
wire open_36;
wire open_37;
wire open_38;
wire open_39;
wire open_40;
wire open_41;
wire open_42;
wire open_43;
wire open_44;
wire open_45;
wire open_46;
wire open_47;
wire open_48;
wire open_49;
wire open_50;
wire open_51;
wire open_52;
wire open_53;
wire open_54;
wire open_55;
wire open_56;
wire open_57;
wire open_58;
wire open_59;
wire open_60;
wire open_61;
wire open_62;
wire open_63;
wire open_64;
wire open_65;
wire open_66;
wire open_67;
wire open_68;
wire open_69;
wire open_70;
wire open_71;
wire open_72;
wire open_73;
wire open_74;
wire open_75;
wire open_76;
wire open_77;
wire open_78;
wire open_79;
wire open_80;
wire open_81;
wire open_82;
wire open_83;
wire open_84;
wire open_85;
wire open_86;
wire open_87;
wire open_88;
wire open_89;
wire open_90;
wire open_91;
wire open_92;
wire open_93;
wire open_94;
wire open_95;
wire open_96;
wire open_97;
wire open_98;
wire open_99;
wire open_100;
wire open_101;
wire open_102;
wire open_103;
wire open_104;
wire open_105;
wire open_106;
wire open_107;
wire open_108;
wire open_109;
wire open_110;
wire open_111;
wire open_112;
wire open_113;
wire open_114;
wire open_115;
wire open_116;
wire open_117;
wire open_118;
wire open_119;
wire open_120;
wire open_121;
wire open_122;
wire open_123;
wire open_124;
wire open_125;
wire open_126;
wire open_127;
wire open_128;
wire open_129;
wire open_130;
wire open_131;
wire open_132;
wire open_133;
wire open_134;
wire open_135;
wire open_136;
wire open_137;
wire open_138;
wire open_139;
wire open_140;
wire open_141;
wire open_142;
wire open_143;
wire open_144;
wire open_145;
wire open_146;
wire open_147;
wire open_148;
wire open_149;
wire open_150;
wire open_151;
wire open_152;
wire open_153;
wire open_154;
wire open_155;
wire open_156;
wire open_157;
wire open_158;
wire open_159;
wire open_160;
wire open_161;
wire open_162;
wire open_163;
wire open_164;
wire open_165;
wire open_166;
wire open_167;
wire open_168;
wire open_169;
wire open_170;
wire open_171;
wire open_172;
wire open_173;
wire open_174;
wire open_175;
wire open_176;
wire open_177;
wire open_178;
wire open_179;
wire open_180;
wire open_181;
wire open_182;
wire open_183;
wire open_184;
wire open_185;
wire open_186;
wire open_187;
wire open_188;
wire open_189;
wire open_190;
wire open_191;
wire open_192;
wire open_193;
wire open_194;
wire open_195;
wire open_196;
wire open_197;
wire open_198;
wire open_199;
wire open_200;
wire open_201;
wire open_202;
wire open_203;
wire open_204;
wire open_205;
wire open_206;
wire open_207;
wire open_208;
wire open_209;
wire open_210;
wire open_211;
wire open_212;
wire open_213;
wire open_214;
wire open_215;
wire open_216;
wire open_217;
wire open_218;
wire open_219;
wire open_220;
wire open_221;
wire open_222;
wire open_223;
wire open_224;
wire open_225;
wire open_226;
wire open_227;
wire open_228;
wire open_229;
wire open_230;
wire open_231;
wire open_232;
wire open_233;
wire open_234;
wire open_235;
wire open_236;
wire open_237;
wire open_238;
wire open_239;
wire n210;
// (18, 11, 'lutff_6/cout')

wire n211;
// (21, 20, 'lutff_5/cout')

wire n212;
// (18, 11, 'lutff_0/cout')

wire n213;
// (18, 12, 'lutff_0/cout')

wire n214;
// (18, 11, 'lutff_2/cout')

wire n215;
// (18, 12, 'lutff_2/cout')

wire n216;
// (18, 12, 'lutff_4/cout')

wire n217;
// (21, 21, 'lutff_0/cout')

wire n218;
// (18, 12, 'lutff_6/cout')

wire n219;
// (21, 19, 'lutff_3/cout')

wire n220;
// (22, 21, 'lutff_0/cout')

wire n221;
// (21, 19, 'lutff_1/cout')

wire n222;
// (22, 19, 'lutff_0/cout')

wire n223;
// (22, 19, 'lutff_2/cout')

wire n224;
// (21, 19, 'lutff_5/cout')

wire n225;
// (22, 19, 'lutff_4/cout')

wire n226;
// (22, 20, 'lutff_5/cout')

wire n227;
// (22, 19, 'lutff_6/cout')

wire n228;
// (7, 20, 'lutff_0/cout')

wire n229;
// (18, 13, 'lutff_0/cout')

wire n230;
// (22, 20, 'lutff_1/cout')

wire n231;
// (22, 20, 'lutff_3/cout')

wire n232;
// (21, 20, 'lutff_2/cout')

wire n233;
// (21, 20, 'lutff_0/cout')

wire n234;
// (21, 20, 'lutff_6/cout')

wire n235;
// (18, 11, 'lutff_5/cout')

wire n236;
// (21, 20, 'lutff_4/cout')

wire n237;
// (18, 12, 'lutff_1/cout')

wire n238;
// (18, 11, 'lutff_1/cout')

wire n239;
// (18, 12, 'lutff_3/cout')

wire n240;
// (18, 11, 'lutff_3/cout')

wire n241;
// (18, 12, 'lutff_5/cout')

wire n242;
// (16, 14, 'lutff_0/cout')

wire n243;
// (16, 11, 'lutff_0/cout')

wire n244;
// (21, 19, 'lutff_2/cout')

wire n245;
// (21, 19, 'lutff_0/cout')

wire n246;
// (22, 19, 'lutff_1/cout')

wire n247;
// (21, 19, 'lutff_6/cout')

wire n248;
// (22, 19, 'lutff_3/cout')

wire n249;
// (21, 19, 'lutff_4/cout')

wire n250;
// (22, 19, 'lutff_5/cout')

wire n251;
// (22, 20, 'lutff_4/cout')

wire n252;
// (22, 20, 'lutff_6/cout')

wire n253;
// (22, 20, 'lutff_0/cout')

wire n254;
// (21, 20, 'lutff_3/cout')

wire n255;
// (22, 20, 'lutff_2/cout')

wire n256;
// (21, 20, 'lutff_1/cout')

wire n257;
// (18, 11, 'lutff_4/cout')

wire n258;
// (18, 11, 'lutff_6/out')

wire n259;
// (18, 11, 'lutff_6/lout')

wire n260;
// (16, 12, 'lutff_4/lout')

wire n261;
// (21, 20, 'lutff_5/out')

wire n262;
// (21, 20, 'lutff_5/lout')

wire n263;
// (7, 21, 'lutff_2/lout')

wire n264;
// (17, 11, 'lutff_1/lout')

wire n265;
// (7, 19, 'lutff_2/lout')

wire n266;
// (18, 11, 'lutff_0/out')

wire n267;
// (18, 11, 'lutff_0/lout')

wire n268;
// (18, 11, 'carry_in_mux')

// Carry-In for (18 11)
assign n268 = 1;

wire n269;
// (24, 22, 'lutff_5/lout')

wire n270;
// (16, 14, 'lutff_5/lout')

wire n271;
// (18, 12, 'lutff_0/out')

wire n272;
// (18, 12, 'lutff_0/lout')

wire n273;
// (18, 11, 'lutff_2/out')

wire n274;
// (18, 11, 'lutff_2/lout')

wire n275;
// (24, 22, 'lutff_7/lout')

wire n276;
// (18, 12, 'lutff_2/out')

wire n277;
// (18, 12, 'lutff_2/lout')

wire n278;
// (9, 25, 'lutff_6/lout')

wire n279;
// (16, 14, 'lutff_1/out')

wire n280;
// (16, 14, 'lutff_1/lout')

wire n281;
// (18, 12, 'lutff_4/out')

wire n282;
// (18, 12, 'lutff_4/lout')

wire n283;
// (16, 11, 'lutff_3/lout')

wire n284;
// (21, 21, 'lutff_0/lout')

wire n285;
// (16, 14, 'lutff_3/lout')

wire n286;
// (18, 12, 'lutff_6/out')

wire n287;
// (18, 12, 'lutff_6/lout')

wire n288;
// (26, 20, 'lutff_6/lout')

wire n289;
// (16, 11, 'lutff_1/out')

wire n290;
// (16, 11, 'lutff_1/lout')

wire n291;
// (22, 21, 'lutff_6/lout')

wire n292;
// (24, 25, 'lutff_5/lout')

wire n293;
// (16, 11, 'lutff_7/lout')

wire n294;
// (23, 20, 'lutff_2/lout')

wire n295;
// (22, 21, 'lutff_4/lout')

wire n296;
// (24, 25, 'lutff_7/lout')

wire n297;
// (19, 12, 'lutff_5/lout')

wire n298;
// (16, 11, 'lutff_5/lout')

wire n299;
// (23, 20, 'lutff_4/lout')

wire n300;
// (18, 10, 'lutff_7/lout')

wire n301;
// (21, 19, 'lutff_3/out')

wire n302;
// (21, 19, 'lutff_3/lout')

wire n303;
// (24, 21, 'lutff_4/lout')

wire n304;
// (9, 19, 'lutff_1/lout')

wire n305;
// (23, 20, 'lutff_6/lout')

wire n306;
// (15, 15, 'lutff_5/lout')

wire n307;
// (7, 23, 'lutff_5/lout')

wire n308;
// (22, 21, 'lutff_0/lout')

wire n309;
// (17, 12, 'lutff_7/lout')

wire n310;
// (18, 10, 'lutff_5/lout')

wire n311;
// (21, 19, 'lutff_1/out')

wire n312;
// (21, 19, 'lutff_1/lout')

wire n313;
// (17, 12, 'lutff_5/lout')

wire n314;
// (22, 19, 'lutff_0/out')

wire n315;
// (22, 19, 'lutff_0/lout')

wire n316;
// (22, 19, 'carry_in_mux')

// Carry-In for (22 19)
assign n316 = 1;

wire n317;
// (22, 22, 'lutff_6/lout')

wire n318;
// (21, 19, 'lutff_7/out')

wire n319;
// (21, 19, 'lutff_7/lout')

wire n320;
// (17, 12, 'lutff_3/lout')

wire n321;
// (22, 19, 'lutff_2/out')

wire n322;
// (22, 19, 'lutff_2/lout')

wire n323;
// (20, 19, 'lutff_7/lout')

wire n324;
// (24, 21, 'lutff_2/lout')

wire n325;
// (21, 19, 'lutff_5/out')

wire n326;
// (21, 19, 'lutff_5/lout')

wire n327;
// (23, 21, 'lutff_1/lout')

wire n328;
// (1, 23, 'lutff_0/lout')

wire n329;
// (17, 12, 'lutff_1/lout')

wire n330;
// (22, 19, 'lutff_4/out')

wire n331;
// (22, 19, 'lutff_4/lout')

wire n332;
// (20, 19, 'lutff_5/lout')

wire n333;
// (22, 20, 'lutff_5/out')

wire n334;
// (22, 20, 'lutff_5/lout')

wire n335;
// (26, 21, 'lutff_2/lout')

wire n336;
// (22, 18, 'lutff_7/lout')

wire n337;
// (22, 19, 'lutff_6/out')

wire n338;
// (22, 19, 'lutff_6/lout')

wire n339;
// (22, 20, 'lutff_7/out')

wire n340;
// (22, 20, 'lutff_7/lout')

wire n341;
// (7, 20, 'lutff_0/out')

wire n342;
// (7, 20, 'lutff_0/lout')

wire n343;
// (7, 20, 'carry_in_mux')

// Carry-In for (7 20)
assign n343 = 1;

wire n344;
// (22, 18, 'lutff_5/lout')

wire n345;
// (18, 13, 'lutff_0/lout')

wire n346;
// (22, 20, 'lutff_1/out')

wire n347;
// (22, 20, 'lutff_1/lout')

wire n348;
// (17, 10, 'lutff_3/lout')

wire n349;
// (7, 20, 'lutff_2/lout')

wire n350;
// (24, 26, 'lutff_1/lout')

wire n351;
// (16, 20, 'lutff_4/lout')

wire n352;
// (16, 12, 'lutff_3/lout')

wire n353;
// (11, 24, 'lutff_7/lout')

wire n354;
// (22, 20, 'lutff_3/out')

wire n355;
// (22, 20, 'lutff_3/lout')

wire n356;
// (16, 15, 'lutff_3/lout')

wire n357;
// (6, 21, 'lutff_2/lout')

wire n358;
// (7, 20, 'lutff_4/lout')

wire n359;
// (21, 20, 'lutff_2/out')

wire n360;
// (21, 20, 'lutff_2/lout')

wire n361;
// (16, 12, 'lutff_1/lout')

wire n362;
// (17, 11, 'lutff_6/lout')

wire n363;
// (7, 21, 'lutff_7/lout')

wire n364;
// (24, 20, 'lutff_1/lout')

wire n365;
// (7, 20, 'lutff_6/lout')

wire n366;
// (21, 20, 'lutff_0/out')

wire n367;
// (21, 20, 'lutff_0/lout')

wire n368;
// (16, 12, 'lutff_7/lout')

wire n369;
// (17, 11, 'lutff_4/lout')

wire n370;
// (7, 21, 'lutff_5/lout')

wire n371;
// (21, 20, 'lutff_6/out')

wire n372;
// (21, 20, 'lutff_6/lout')

wire n373;
// (17, 13, 'lutff_0/lout')

wire n374;
// (18, 11, 'lutff_5/out')

wire n375;
// (18, 11, 'lutff_5/lout')

wire n376;
// (16, 12, 'lutff_5/lout')

wire n377;
// (17, 11, 'lutff_2/lout')

wire n378;
// (21, 20, 'lutff_4/out')

wire n379;
// (21, 20, 'lutff_4/lout')

wire n380;
// (9, 23, 'lutff_3/lout')

wire n381;
// (7, 19, 'lutff_3/lout')

wire n382;
// (26, 19, 'lutff_7/lout')

wire n383;
// (18, 11, 'lutff_7/out')

wire n384;
// (18, 11, 'lutff_7/lout')

wire n385;
// (17, 11, 'lutff_0/lout')

wire n386;
// (7, 21, 'lutff_1/lout')

wire n387;
// (7, 22, 'lutff_1/lout')

wire n388;
// (18, 12, 'lutff_1/out')

wire n389;
// (18, 12, 'lutff_1/lout')

wire n390;
// (24, 17, 'lutff_5/lout')

wire n391;
// (18, 11, 'lutff_1/out')

wire n392;
// (18, 11, 'lutff_1/lout')

wire n393;
// (16, 14, 'lutff_4/lout')

wire n394;
// (20, 20, 'lutff_2/lout')

wire n395;
// (18, 12, 'lutff_3/out')

wire n396;
// (18, 12, 'lutff_3/lout')

wire n397;
// (24, 17, 'lutff_7/lout')

wire n398;
// (18, 11, 'lutff_3/out')

wire n399;
// (18, 11, 'lutff_3/lout')

wire n400;
// (7, 22, 'lutff_5/lout')

wire n401;
// (18, 12, 'lutff_5/out')

wire n402;
// (18, 12, 'lutff_5/lout')

wire n403;
// (16, 11, 'lutff_2/lout')

wire n404;
// (16, 14, 'lutff_0/out')

wire n405;
// (16, 14, 'lutff_0/lout')

wire n406;
// (16, 14, 'carry_in_mux')

// Carry-In for (16 14)
assign n406 = 1;

wire n407;
// (6, 20, 'lutff_1/lout')

wire n408;
// (18, 12, 'lutff_7/out')

wire n409;
// (18, 12, 'lutff_7/lout')

wire n410;
// (16, 11, 'lutff_0/out')

wire n411;
// (16, 11, 'lutff_0/lout')

wire n412;
// (16, 11, 'carry_in_mux')

// Carry-In for (16 11)
assign n412 = 1;

wire n413;
// (21, 18, 'lutff_3/lout')

wire n414;
// (16, 14, 'lutff_2/lout')

wire n415;
// (16, 11, 'lutff_6/lout')

wire n416;
// (18, 10, 'lutff_2/lout')

wire n417;
// (16, 11, 'lutff_4/lout')

wire n418;
// (22, 21, 'lutff_5/lout')

wire n419;
// (7, 23, 'lutff_0/lout')

wire n420;
// (18, 10, 'lutff_0/lout')

wire n421;
// (18, 23, 'lutff_7/lout')

wire n422;
// (22, 21, 'lutff_3/lout')

wire n423;
// (9, 19, 'lutff_2/lout')

wire n424;
// (17, 12, 'lutff_6/lout')

wire n425;
// (7, 25, 'lutff_0/lout')

wire n426;
// (23, 21, 'lutff_6/lout')

wire n427;
// (16, 13, 'lutff_5/lout')

wire n428;
// (9, 19, 'lutff_0/lout')

wire n429;
// (21, 19, 'lutff_2/out')

wire n430;
// (21, 19, 'lutff_2/lout')

wire n431;
// (15, 15, 'lutff_4/lout')

wire n432;
// (17, 12, 'lutff_4/lout')

wire n433;
// (18, 10, 'lutff_4/lout')

wire n434;
// (24, 21, 'lutff_7/lout')

wire n435;
// (21, 19, 'lutff_0/out')

wire n436;
// (21, 19, 'lutff_0/lout')

wire n437;
// (21, 19, 'carry_in_mux')

// Carry-In for (21 19)
assign n437 = 1;

wire n438;
// (7, 23, 'lutff_6/lout')

wire n439;
// (17, 12, 'lutff_2/lout')

wire n440;
// (22, 19, 'lutff_1/out')

wire n441;
// (22, 19, 'lutff_1/lout')

wire n442;
// (20, 19, 'lutff_6/lout')

wire n443;
// (21, 19, 'lutff_6/out')

wire n444;
// (21, 19, 'lutff_6/lout')

wire n445;
// (17, 12, 'lutff_0/lout')

wire n446;
// (22, 19, 'lutff_3/out')

wire n447;
// (22, 19, 'lutff_3/lout')

wire n448;
// (17, 21, 'lutff_4/lout')

wire n449;
// (23, 21, 'lutff_0/lout')

wire n450;
// (21, 19, 'lutff_4/out')

wire n451;
// (21, 19, 'lutff_4/lout')

wire n452;
// (24, 21, 'lutff_3/lout')

wire n453;
// (22, 19, 'lutff_5/out')

wire n454;
// (22, 19, 'lutff_5/lout')

wire n455;
// (22, 20, 'lutff_4/out')

wire n456;
// (22, 20, 'lutff_4/lout')

wire n457;
// (22, 19, 'lutff_7/out')

wire n458;
// (22, 19, 'lutff_7/lout')

wire n459;
// (22, 20, 'lutff_6/out')

wire n460;
// (22, 20, 'lutff_6/lout')

wire n461;
// (17, 10, 'lutff_2/lout')

wire n462;
// (7, 20, 'lutff_1/out')

wire n463;
// (7, 20, 'lutff_1/lout')

wire n464;
// (22, 20, 'lutff_0/out')

wire n465;
// (22, 20, 'lutff_0/lout')

wire n466;
// (16, 15, 'lutff_2/lout')

wire n467;
// (7, 20, 'lutff_3/lout')

wire n468;
// (30, 1, 'lutff_6/lout')

wire n469;
// (24, 26, 'lutff_0/lout')

wire n470;
// (17, 13, 'lutff_5/lout')

wire n471;
// (22, 18, 'lutff_2/lout')

wire n472;
// (16, 12, 'lutff_2/lout')

wire n473;
// (17, 11, 'lutff_7/lout')

wire n474;
// (21, 20, 'lutff_3/out')

wire n475;
// (21, 20, 'lutff_3/lout')

wire n476;
// (22, 20, 'lutff_2/out')

wire n477;
// (22, 20, 'lutff_2/lout')

wire n478;
// (6, 21, 'lutff_3/lout')

wire n479;
// (7, 20, 'lutff_5/lout')

wire n480;
// (17, 13, 'lutff_7/lout')

wire n481;
// (7, 19, 'lutff_4/lout')

wire n482;
// (22, 18, 'lutff_0/lout')

wire n483;
// (16, 12, 'lutff_0/lout')

wire n484;
// (12, 23, 'lutff_0/lout')

wire n485;
// (7, 21, 'lutff_6/lout')

wire n486;
// (17, 11, 'lutff_5/lout')

wire n487;
// (7, 20, 'lutff_7/lout')

wire n488;
// (21, 20, 'lutff_1/out')

wire n489;
// (21, 20, 'lutff_1/lout')

wire n490;
// (18, 11, 'lutff_4/out')

wire n491;
// (18, 11, 'lutff_4/lout')

wire n492;
// (16, 12, 'lutff_6/lout')

wire n493;
// (17, 11, 'lutff_3/lout')

wire n494;
// (7, 21, 'lutff_4/lout')

wire n495;
// (21, 20, 'lutff_7/out')

wire n496;
// (21, 20, 'lutff_7/lout')

wire n497;
// (24, 20, 'lutff_6/lout')

wire n498;
// (17, 13, 'lutff_3/lout')

wire n499;
// (7, 19, 'lutff_0/lout')

// RAM TILE 8 15
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_15 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_0, open_1, open_2, open_3, n53, open_4, open_5, open_6, open_7, open_8, open_9, open_10, n54, open_12, open_13, open_14}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n52),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 15
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_15 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_15, open_16, open_17, open_18, n193, open_19, open_20, open_21, open_22, open_23, open_24, open_25, n194, open_27, open_28, open_29}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n52),
  .RCLK(io_0_27_1)
);

// RAM TILE 8 17
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_17 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_30, open_31, open_32, open_33, n56, open_34, open_35, open_36, open_37, open_38, open_39, open_40, n57, open_42, open_43, open_44}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n66),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 17
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000101000100000100),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_17 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_45, open_46, open_47, open_48, n195, open_49, open_50, open_51, open_52, open_53, open_54, open_55, n196, open_57, open_58, open_59}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n189),
  .RCLK(io_0_27_1)
);

// RAM TILE 8 19
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_19 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_60, open_61, open_62, open_63, n60, open_64, open_65, open_66, open_67, open_68, open_69, open_70, n64, open_72, open_73, open_74}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n59),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 19
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000010000000101),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_19 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, n208, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_75, open_76, open_77, open_78, n28, open_79, open_80, open_81, open_82, open_83, open_84, open_85, n87, open_87, open_88, open_89}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n189),
  .RCLK(io_0_27_1)
);

// RAM TILE 8 21
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_21 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_90, open_91, open_92, open_93, n73, open_94, open_95, open_96, open_97, open_98, open_99, open_100, n74, open_102, open_103, open_104}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n66),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 21
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_21 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_105, open_106, open_107, open_108, n197, open_109, open_110, open_111, open_112, open_113, open_114, open_115, n200, open_117, open_118, open_119}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n52),
  .RCLK(io_0_27_1)
);

// RAM TILE 8 23
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_23 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_120, open_121, open_122, open_123, n76, open_124, open_125, open_126, open_127, open_128, open_129, open_130, n78, open_132, open_133, open_134}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n66),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 23
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000100000100),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_23 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_135, open_136, open_137, open_138, n198, open_139, open_140, open_141, open_142, open_143, open_144, open_145, n201, open_147, open_148, open_149}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n189),
  .RCLK(io_0_27_1)
);

// RAM TILE 8 25
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_25 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_150, open_151, open_152, open_153, n81, open_154, open_155, open_156, open_157, open_158, open_159, open_160, n83, open_162, open_163, open_164}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n66),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 25
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_25 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_165, open_166, open_167, open_168, n203, open_169, open_170, open_171, open_172, open_173, open_174, open_175, n204, open_177, open_178, open_179}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n52),
  .RCLK(io_0_27_1)
);

// RAM TILE 8 27
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_27 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_180, open_181, open_182, open_183, n82, open_184, open_185, open_186, open_187, open_188, open_189, open_190, n84, open_192, open_193, open_194}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n59),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 27
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000101000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_27 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_195, open_196, open_197, open_198, n206, open_199, open_200, open_201, open_202, open_203, open_204, open_205, n205, open_207, open_208, open_209}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n189),
  .RCLK(io_0_27_1)
);

// RAM TILE 8 29
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_8_29 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_210, open_211, open_212, open_213, n77, open_214, open_215, open_216, open_217, open_218, open_219, open_220, n79, open_222, open_223, open_224}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n59),
  .RCLK(io_0_27_1)
);

// RAM TILE 25 29
SB_RAM40_4K #(
  .READ_MODE(3),
  .WRITE_MODE(3),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_25_29 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RADDR({io_33_27_1, io_33_30_0, io_33_29_1, io_33_31_0, io_33_30_1, io_31_33_0, io_31_33_1, io_30_33_0, io_30_33_1, io_4_33_0, io_3_33_1}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({open_225, open_226, open_227, open_228, n207, open_229, open_230, open_231, open_232, open_233, open_234, open_235, n202, open_237, open_238, open_239}),
  .WE(io_0_11_0),
  .WCLKE(io_0_16_0),
  .WCLK(io_0_16_0),
  .RE(io_0_11_0),
  .RCLKE(n59),
  .RCLK(io_0_27_1)
);

assign n259 = /* LUT   18 11  6 */ 1'b0;
assign n262 = /* LUT   21 20  5 */ 1'b0;
assign n267 = /* LUT   18 11  0 */ 1'b0;
assign n272 = /* LUT   18 12  0 */ 1'b0;
assign n274 = /* LUT   18 11  2 */ 1'b0;
assign n277 = /* LUT   18 12  2 */ 1'b0;
assign n280 = /* LUT   16 14  1 */ 1'b0;
assign n282 = /* LUT   18 12  4 */ 1'b0;
assign n287 = /* LUT   18 12  6 */ 1'b0;
assign n290 = /* LUT   16 11  1 */ 1'b0;
assign n302 = /* LUT   21 19  3 */ 1'b0;
assign n312 = /* LUT   21 19  1 */ 1'b0;
assign n315 = /* LUT   22 19  0 */ 1'b0;
assign n319 = /* LUT   21 19  7 */ 1'b0;
assign n322 = /* LUT   22 19  2 */ 1'b0;
assign n326 = /* LUT   21 19  5 */ 1'b0;
assign n331 = /* LUT   22 19  4 */ 1'b0;
assign n334 = /* LUT   22 20  5 */ 1'b0;
assign n338 = /* LUT   22 19  6 */ 1'b0;
assign n340 = /* LUT   22 20  7 */ 1'b0;
assign n342 = /* LUT    7 20  0 */ 1'b0;
assign n347 = /* LUT   22 20  1 */ 1'b0;
assign n355 = /* LUT   22 20  3 */ 1'b0;
assign n360 = /* LUT   21 20  2 */ 1'b0;
assign n367 = /* LUT   21 20  0 */ 1'b0;
assign n372 = /* LUT   21 20  6 */ 1'b0;
assign n375 = /* LUT   18 11  5 */ 1'b0;
assign n379 = /* LUT   21 20  4 */ 1'b0;
assign n384 = /* LUT   18 11  7 */ 1'b0;
assign n389 = /* LUT   18 12  1 */ 1'b0;
assign n392 = /* LUT   18 11  1 */ 1'b0;
assign n396 = /* LUT   18 12  3 */ 1'b0;
assign n399 = /* LUT   18 11  3 */ 1'b0;
assign n402 = /* LUT   18 12  5 */ 1'b0;
assign n405 = /* LUT   16 14  0 */ 1'b0;
assign n409 = /* LUT   18 12  7 */ 1'b0;
assign n411 = /* LUT   16 11  0 */ 1'b0;
assign n430 = /* LUT   21 19  2 */ 1'b0;
assign n436 = /* LUT   21 19  0 */ 1'b0;
assign n441 = /* LUT   22 19  1 */ 1'b0;
assign n444 = /* LUT   21 19  6 */ 1'b0;
assign n447 = /* LUT   22 19  3 */ 1'b0;
assign n451 = /* LUT   21 19  4 */ 1'b0;
assign n454 = /* LUT   22 19  5 */ 1'b0;
assign n456 = /* LUT   22 20  4 */ 1'b0;
assign n458 = /* LUT   22 19  7 */ 1'b0;
assign n460 = /* LUT   22 20  6 */ 1'b0;
assign n463 = /* LUT    7 20  1 */ 1'b0;
assign n465 = /* LUT   22 20  0 */ 1'b0;
assign n475 = /* LUT   21 20  3 */ 1'b0;
assign n477 = /* LUT   22 20  2 */ 1'b0;
assign n484 = /* LUT   12 23  0 */ 1'b0;
assign n489 = /* LUT   21 20  1 */ 1'b0;
assign n491 = /* LUT   18 11  4 */ 1'b0;
assign n496 = /* LUT   21 20  7 */ 1'b0;
assign n260 = /* LUT   16 12  4 */ (n139 ? (n101 ? io_0_11_0 : !io_0_11_0) : (n101 ? !io_0_11_0 : io_0_11_0));
assign n263 = /* LUT    7 21  2 */ (n74 ? n30 : 1'b0);
assign n264 = /* LUT   17 11  1 */ !n94;
assign n265 = /* LUT    7 19  2 */ (n56 ? (n60 ? (n58 ? 1'b0 : !n30) : !n30) : (n60 ? !n58 : 1'b1));
assign n269 = /* LUT   24 22  5 */ n189;
assign n270 = /* LUT   16 14  5 */ (n106 ? (n110 ? (n107 ? !n108 : 1'b0) : 1'b0) : 1'b0);
assign n275 = /* LUT   24 22  7 */ (n80 ? (n201 ? (n200 ? 1'b0 : !n86) : !n200) : (n201 ? !n86 : 1'b1));
assign n278 = /* LUT    9 25  6 */ (n84 ? (n83 ? (n58 ? 1'b0 : !n30) : !n58) : (n83 ? !n30 : 1'b1));
assign n283 = /* LUT   16 11  3 */ (n123 ? (io_0_11_0 ? n92 : !n92) : (io_0_11_0 ? !n92 : n92));
assign n284 = /* LUT   21 21  0 */ n176;
assign n285 = /* LUT   16 14  3 */ (n107 ? !io_0_11_0 : io_0_11_0);
assign n288 = /* LUT   26 20  6 */ !io_33_21_1;
assign n291 = /* LUT   22 21  6 */ !io_33_23_1;
assign n292 = /* LUT   24 25  5 */ (n204 ? (n191 ? !n80 : 1'b0) : n191);
assign n293 = /* LUT   16 11  7 */ (n127 ? (io_0_11_0 ? n96 : !n96) : (io_0_11_0 ? !n96 : n96));
assign n294 = /* LUT   23 20  2 */ (io_33_21_1 ? !io_33_28_0 : 1'b0);
assign n295 = /* LUT   22 21  4 */ (n179 ? (io_33_23_1 ? (n184 ? 1'b0 : !n177) : (n184 ? 1'b1 : !n177)) : !n177);
assign n296 = /* LUT   24 25  7 */ (n192 ? (n80 ? !n203 : 1'b1) : 1'b0);
assign n297 = /* LUT   19 12  5 */ !n154;
assign n298 = /* LUT   16 11  5 */ (n125 ? (n94 ? io_0_11_0 : !io_0_11_0) : (n94 ? !io_0_11_0 : io_0_11_0));
assign n299 = /* LUT   23 20  4 */ (io_33_28_0 ? io_33_21_1 : 1'b0);
assign n300 = /* LUT   18 10  7 */ (n154 ? n1 : !n119);
assign n303 = /* LUT   24 21  4 */ (io_33_28_0 ? 1'b0 : !io_33_21_1);
assign n304 = /* LUT    9 19  1 */ (n54 ? (n85 ? !n80 : 1'b0) : n85);
assign n305 = /* LUT   23 20  6 */ !io_33_28_0;
assign n306 = /* LUT   15 15  5 */ io_0_27_1;
assign n307 = /* LUT    7 23  5 */ (n75 ? (n79 ? !n58 : 1'b1) : 1'b0);
assign n308 = /* LUT   22 21  0 */ n182;
assign n309 = /* LUT   17 12  7 */ !n103;
assign n310 = /* LUT   18 10  5 */ !n105;
assign n313 = /* LUT   17 12  5 */ (n102 ? 1'b0 : (n104 ? 1'b0 : (n103 ? 1'b0 : !n101)));
assign n317 = /* LUT   22 22  6 */ io_33_30_1;
assign n320 = /* LUT   17 12  3 */ (n1 ? 1'b1 : !n154);
assign n323 = /* LUT   20 19  7 */ !io_31_33_0;
assign n324 = /* LUT   24 21  2 */ (io_33_20_1 ? 1'b0 : (io_33_21_0 ? 1'b0 : (io_33_27_1 ? 1'b0 : n190)));
assign n327 = /* LUT   23 21  1 */ (n185 ? n183 : 1'b0);
assign n328 = /* LUT    1 23  0 */ (io_0_27_0 ? (io_0_11_1 ? 1'b0 : io_0_25_0) : 1'b0);
assign n329 = /* LUT   17 12  1 */ !n100;
assign n332 = /* LUT   20 19  5 */ !io_33_31_0;
assign n335 = /* LUT   26 21  2 */ (io_33_30_0 ? 1'b0 : (io_33_28_0 ? 1'b0 : (io_33_21_1 ? 1'b0 : !io_33_29_1)));
assign n336 = /* LUT   22 18  7 */ !io_3_33_1;
assign n344 = /* LUT   22 18  5 */ !io_33_30_1;
assign n345 = /* LUT   18 13  0 */ n158;
assign n348 = /* LUT   17 10  3 */ !n93;
assign n349 = /* LUT    7 20  2 */ (n67 ? !n38 : n38);
assign n350 = /* LUT   24 26  1 */ (n207 ? (n86 ? (n58 ? 1'b0 : !n206) : !n58) : (n86 ? !n206 : 1'b1));
assign n351 = /* LUT   16 20  4 */ n59;
assign n352 = /* LUT   16 12  3 */ (n138 ? (io_0_11_0 ? n100 : !n100) : (io_0_11_0 ? !n100 : n100));
assign n353 = /* LUT   11 24  7 */ 1'b1;
assign n356 = /* LUT   16 15  3 */ !n110;
assign n357 = /* LUT    6 21  2 */ (n18 ? n27 : 1'b0);
assign n358 = /* LUT    7 20  4 */ (n69 ? !n40 : n40);
assign n361 = /* LUT   16 12  1 */ (n136 ? (io_0_11_0 ? n98 : !n98) : (io_0_11_0 ? !n98 : n98));
assign n362 = /* LUT   17 11  6 */ (n131 ? (io_29_0_0 ? (n120 ? n153 : 1'b0) : 1'b1) : 1'b0);
assign n363 = /* LUT    7 21  7 */ (n42 ? (n61 ? (n44 ? 1'b1 : n18) : 1'b1) : (n61 ? (n44 ? !n18 : 1'b0) : !n18));
assign n364 = /* LUT   24 20  1 */ (io_33_21_1 ? 1'b0 : io_33_28_0);
assign n365 = /* LUT    7 20  6 */ (n71 ? !n42 : n42);
assign n368 = /* LUT   16 12  7 */ (n142 ? (n104 ? io_0_11_0 : !io_0_11_0) : (n104 ? !io_0_11_0 : io_0_11_0));
assign n369 = /* LUT   17 11  4 */ !n92;
assign n370 = /* LUT    7 21  5 */ (n43 ? (n18 ? 1'b1 : (n45 ? 1'b1 : !n65)) : (n18 ? 1'b0 : (n45 ? 1'b1 : !n65)));
assign n373 = /* LUT   17 13  0 */ !n99;
assign n376 = /* LUT   16 12  5 */ (n140 ? (io_0_11_0 ? n102 : !n102) : (io_0_11_0 ? !n102 : n102));
assign n377 = /* LUT   17 11  2 */ (n96 ? 1'b0 : (n93 ? 1'b0 : (n94 ? 1'b0 : !n95)));
assign n380 = /* LUT    9 23  3 */ (n80 ? 1'b0 : (n86 ? 1'b0 : !n58));
assign n381 = /* LUT    7 19  3 */ (n41 ? (n37 ? (n18 ? 1'b1 : !n62) : 1'b1) : (n37 ? (n18 ? 1'b0 : !n62) : !n18));
assign n382 = /* LUT   26 19  7 */ io_33_30_1;
assign n385 = /* LUT   17 11  0 */ !n95;
assign n386 = /* LUT    7 21  1 */ (n32 ? (n25 ? (n46 ? n18 : 1'b1) : 1'b1) : (n25 ? (n46 ? 1'b0 : !n18) : !n18));
assign n387 = /* LUT    7 22  1 */ (n18 ? n27 : !n49);
assign n390 = /* LUT   24 17  5 */ (n195 ? (n193 ? (n86 ? 1'b0 : !n80) : !n86) : (n193 ? !n80 : 1'b1));
assign n393 = /* LUT   16 14  4 */ (n89 ? n4 : !n4);
assign n394 = /* LUT   20 20  2 */ !io_33_30_0;
assign n397 = /* LUT   24 17  7 */ (n194 ? (n80 ? 1'b0 : (n86 ? !n196 : 1'b1)) : (n86 ? !n196 : 1'b1));
assign n400 = /* LUT    7 22  5 */ (n33 ? (n38 ? (n22 ? n18 : 1'b1) : (n22 ? 1'b0 : !n18)) : (n38 ? 1'b1 : !n18));
assign n403 = /* LUT   16 11  2 */ (n122 ? (io_0_11_0 ? n91 : !n91) : (io_0_11_0 ? !n91 : n91));
assign n407 = /* LUT    6 20  1 */ (io_0_11_0 ? !n27 : n27);
assign n413 = /* LUT   21 18  3 */ !io_4_33_0;
assign n414 = /* LUT   16 14  2 */ (n147 ? !n106 : n106);
assign n415 = /* LUT   16 11  6 */ (n126 ? (io_0_11_0 ? n95 : !n95) : (io_0_11_0 ? !n95 : n95));
assign n416 = /* LUT   18 10  2 */ n152;
assign n417 = /* LUT   16 11  4 */ (n124 ? (io_0_11_0 ? n93 : !n93) : (io_0_11_0 ? !n93 : n93));
assign n418 = /* LUT   22 21  5 */ !io_33_29_1;
assign n419 = /* LUT    7 23  0 */ (n30 ? (n58 ? (n77 ? 1'b0 : !n76) : !n76) : (n58 ? !n77 : 1'b1));
assign n420 = /* LUT   18 10  0 */ !n119;
assign n421 = /* LUT   18 23  7 */ n52;
assign n422 = /* LUT   22 21  3 */ !io_33_27_1;
assign n423 = /* LUT    9 19  2 */ (n87 ? (n86 ? 1'b0 : (n58 ? !n64 : 1'b1)) : (n58 ? !n64 : 1'b1));
assign n424 = /* LUT   17 12  6 */ (n99 ? 1'b0 : (n98 ? 1'b0 : (n100 ? 1'b0 : !n97)));
assign n425 = /* LUT    7 25  0 */ (n81 ? (n30 ? 1'b0 : (n58 ? !n82 : 1'b1)) : (n58 ? !n82 : 1'b1));
assign n426 = /* LUT   23 21  6 */ (io_30_33_0 ? 1'b0 : (io_3_33_1 ? 1'b0 : (io_30_33_1 ? 1'b0 : !io_4_33_0)));
assign n427 = /* LUT   16 13  5 */ !n4;
assign n428 = /* LUT    9 19  0 */ (n80 ? (n86 ? (n53 ? 1'b0 : !n28) : !n53) : (n86 ? !n28 : 1'b1));
assign n431 = /* LUT   15 15  4 */ n90;
assign n432 = /* LUT   17 12  4 */ !n101;
assign n433 = /* LUT   18 10  4 */ n151;
assign n434 = /* LUT   24 21  7 */ (n86 ? (n197 ? (n80 ? 1'b0 : !n198) : !n198) : (n197 ? !n80 : 1'b1));
assign n438 = /* LUT    7 23  6 */ (n48 ? (n30 ? !n78 : 1'b1) : 1'b0);
assign n439 = /* LUT   17 12  2 */ (n134 ? (n116 ? (n133 ? n115 : 1'b0) : 1'b0) : 1'b0);
assign n442 = /* LUT   20 19  6 */ !io_31_33_1;
assign n445 = /* LUT   17 12  0 */ !n102;
assign n448 = /* LUT   17 21  4 */ (io_0_27_0 ? 1'b0 : n155);
assign n449 = /* LUT   23 21  0 */ (io_31_33_0 ? 1'b0 : (io_33_31_0 ? 1'b0 : (io_31_33_1 ? 1'b0 : !n178)));
assign n452 = /* LUT   24 21  3 */ !io_33_21_0;
assign n461 = /* LUT   17 10  2 */ !n91;
assign n466 = /* LUT   16 15  2 */ (n107 ? 1'b1 : n108);
assign n467 = /* LUT    7 20  3 */ (n68 ? !n39 : n39);
assign n468 = /* LUT   30  1  6 */ n157;
assign n469 = /* LUT   24 26  0 */ (n202 ? (n58 ? 1'b0 : (n86 ? !n205 : 1'b1)) : (n86 ? !n205 : 1'b1));
assign n470 = /* LUT   17 13  5 */ !n104;
assign n471 = /* LUT   22 18  2 */ !io_30_33_0;
assign n472 = /* LUT   16 12  2 */ (n137 ? (io_0_11_0 ? n99 : !n99) : (io_0_11_0 ? !n99 : n99));
assign n473 = /* LUT   17 11  7 */ (n119 ? !io_0_11_0 : io_0_11_0);
assign n478 = /* LUT    6 21  3 */ !n32;
assign n479 = /* LUT    7 20  5 */ (n70 ? !n41 : n41);
assign n480 = /* LUT   17 13  7 */ !n97;
assign n481 = /* LUT    7 19  4 */ (n30 ? n57 : 1'b0);
assign n482 = /* LUT   22 18  0 */ !io_30_33_1;
assign n483 = /* LUT   16 12  0 */ (n128 ? (n97 ? io_0_11_0 : !io_0_11_0) : (n97 ? !io_0_11_0 : io_0_11_0));
assign n485 = /* LUT    7 21  6 */ (n30 ? n73 : 1'b0);
assign n486 = /* LUT   17 11  5 */ !n96;
assign n487 = /* LUT    7 20  7 */ (n72 ? !n43 : n43);
assign n492 = /* LUT   16 12  6 */ (n141 ? (io_0_11_0 ? n103 : !n103) : (io_0_11_0 ? !n103 : n103));
assign n493 = /* LUT   17 11  3 */ (n119 ? 1'b0 : (n105 ? 1'b0 : (n91 ? 1'b0 : !n92)));
assign n494 = /* LUT    7 21  4 */ (n39 ? (n18 ? 1'b1 : (n21 ? !n50 : 1'b1)) : (n18 ? 1'b0 : (n21 ? !n50 : 1'b1)));
assign n497 = /* LUT   24 20  6 */ !io_33_20_1;
assign n498 = /* LUT   17 13  3 */ !n98;
assign n499 = /* LUT    7 19  0 */ (n63 ? (n18 ? n40 : n36) : (n18 ? n40 : 1'b1));
assign n210 = /* CARRY 18 11  6 */ (n113 & 1'b0) | ((n113 | 1'b0) & n235);
assign n140 = /* CARRY 16 12  4 */ (io_0_11_0 & n101) | ((io_0_11_0 | n101) & n139);
assign n211 = /* CARRY 21 20  5 */ (n174 & io_0_11_0) | ((n174 | io_0_11_0) & n236);
assign n212 = /* CARRY 18 11  0 */ (1'b0 & n149) | ((1'b0 | n149) & n268);
assign n213 = /* CARRY 18 12  0 */ (1'b0 & n146) | ((1'b0 | n146) & n156);
assign n214 = /* CARRY 18 11  2 */ (1'b0 & n111) | ((1'b0 | n111) & n238);
assign n215 = /* CARRY 18 12  2 */ (1'b0 & n143) | ((1'b0 | n143) & n237);
assign n147 = /* CARRY 16 14  1 */ (1'b0 & n110) | ((1'b0 | n110) & n242);
assign n216 = /* CARRY 18 12  4 */ (1'b0 & n132) | ((1'b0 | n132) & n239);
assign n124 = /* CARRY 16 11  3 */ (n92 & io_0_11_0) | ((n92 | io_0_11_0) & n123);
assign n217 = /* CARRY 21 21  0 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n176);
assign n218 = /* CARRY 18 12  6 */ (n135 & 1'b0) | ((n135 | 1'b0) & n241);
assign n122 = /* CARRY 16 11  1 */ (io_0_11_0 & n105) | ((io_0_11_0 | n105) & n243);
assign n128 = /* CARRY 16 11  7 */ (n96 & io_0_11_0) | ((n96 | io_0_11_0) & n127);
assign n126 = /* CARRY 16 11  5 */ (io_0_11_0 & n94) | ((io_0_11_0 | n94) & n125);
assign n219 = /* CARRY 21 19  3 */ (1'b0 & n167) | ((1'b0 | n167) & n244);
assign n220 = /* CARRY 22 21  0 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n182);
assign n221 = /* CARRY 21 19  1 */ (n163 & 1'b0) | ((n163 | 1'b0) & n245);
assign n222 = /* CARRY 22 19  0 */ (n169 & 1'b0) | ((n169 | 1'b0) & n316);
assign n170 = /* CARRY 21 19  7 */ (n159 & 1'b0) | ((n159 | 1'b0) & n247);
assign n223 = /* CARRY 22 19  2 */ (1'b0 & n166) | ((1'b0 | n166) & n246);
assign n224 = /* CARRY 21 19  5 */ (n161 & 1'b0) | ((n161 | 1'b0) & n249);
assign n225 = /* CARRY 22 19  4 */ (1'b0 & n160) | ((1'b0 | n160) & n248);
assign n226 = /* CARRY 22 20  5 */ (n174 & 1'b0) | ((n174 | 1'b0) & n251);
assign n227 = /* CARRY 22 19  6 */ (1'b0 & n168) | ((1'b0 | n168) & n250);
assign n182 = /* CARRY 22 20  7 */ (n164 & 1'b0) | ((n164 | 1'b0) & n252);
assign n228 = /* CARRY  7 20  0 */ (1'b0 & n27) | ((1'b0 | n27) & n343);
assign n229 = /* CARRY 18 13  0 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n158);
assign n230 = /* CARRY 22 20  1 */ (n162 & 1'b0) | ((n162 | 1'b0) & n253);
assign n68  = /* CARRY  7 20  2 */ (1'b0 & n38) | ((1'b0 | n38) & n67);
assign n139 = /* CARRY 16 12  3 */ (n100 & io_0_11_0) | ((n100 | io_0_11_0) & n138);
assign n231 = /* CARRY 22 20  3 */ (1'b0 & n172) | ((1'b0 | n172) & n255);
assign n70  = /* CARRY  7 20  4 */ (1'b0 & n40) | ((1'b0 | n40) & n69);
assign n232 = /* CARRY 21 20  2 */ (n173 & 1'b0) | ((n173 | 1'b0) & n256);
assign n137 = /* CARRY 16 12  1 */ (n98 & io_0_11_0) | ((n98 | io_0_11_0) & n136);
assign n72  = /* CARRY  7 20  6 */ (n42 & 1'b0) | ((n42 | 1'b0) & n71);
assign n233 = /* CARRY 21 20  0 */ (1'b0 & n175) | ((1'b0 | n175) & n170);
assign n234 = /* CARRY 21 20  6 */ (n171 & 1'b0) | ((n171 | 1'b0) & n211);
assign n235 = /* CARRY 18 11  5 */ (n114 & 1'b0) | ((n114 | 1'b0) & n257);
assign n141 = /* CARRY 16 12  5 */ (n102 & io_0_11_0) | ((n102 | io_0_11_0) & n140);
assign n236 = /* CARRY 21 20  4 */ (n165 & 1'b0) | ((n165 | 1'b0) & n254);
assign n156 = /* CARRY 18 11  7 */ (n118 & 1'b0) | ((n118 | 1'b0) & n210);
assign n237 = /* CARRY 18 12  1 */ (1'b0 & n144) | ((1'b0 | n144) & n213);
assign n238 = /* CARRY 18 11  1 */ (1'b0 & n151) | ((1'b0 | n151) & n212);
assign n239 = /* CARRY 18 12  3 */ (n130 & 1'b0) | ((n130 | 1'b0) & n215);
assign n240 = /* CARRY 18 11  3 */ (n117 & 1'b0) | ((n117 | 1'b0) & n214);
assign n241 = /* CARRY 18 12  5 */ (1'b0 & n129) | ((1'b0 | n129) & n216);
assign n123 = /* CARRY 16 11  2 */ (n91 & io_0_11_0) | ((n91 | io_0_11_0) & n122);
assign n242 = /* CARRY 16 14  0 */ (1'b0 & n107) | ((1'b0 | n107) & n406);
assign n158 = /* CARRY 18 12  7 */ (1'b0 & n145) | ((1'b0 | n145) & n218);
assign n243 = /* CARRY 16 11  0 */ (1'b0 & n119) | ((1'b0 | n119) & n412);
assign n127 = /* CARRY 16 11  6 */ (n95 & io_0_11_0) | ((n95 | io_0_11_0) & n126);
assign n125 = /* CARRY 16 11  4 */ (n93 & io_0_11_0) | ((n93 | io_0_11_0) & n124);
assign n244 = /* CARRY 21 19  2 */ (1'b0 & n166) | ((1'b0 | n166) & n221);
assign n245 = /* CARRY 21 19  0 */ (n169 & 1'b0) | ((n169 | 1'b0) & n437);
assign n246 = /* CARRY 22 19  1 */ (n163 & 1'b0) | ((n163 | 1'b0) & n222);
assign n247 = /* CARRY 21 19  6 */ (n168 & 1'b0) | ((n168 | 1'b0) & n224);
assign n248 = /* CARRY 22 19  3 */ (1'b0 & n167) | ((1'b0 | n167) & n223);
assign n249 = /* CARRY 21 19  4 */ (n160 & 1'b0) | ((n160 | 1'b0) & n219);
assign n250 = /* CARRY 22 19  5 */ (n161 & 1'b0) | ((n161 | 1'b0) & n225);
assign n251 = /* CARRY 22 20  4 */ (n165 & 1'b0) | ((n165 | 1'b0) & n231);
assign n181 = /* CARRY 22 19  7 */ (1'b0 & n159) | ((1'b0 | n159) & n227);
assign n252 = /* CARRY 22 20  6 */ (1'b0 & n171) | ((1'b0 | n171) & n226);
assign n67  = /* CARRY  7 20  1 */ (n32 & 1'b0) | ((n32 | 1'b0) & n228);
assign n253 = /* CARRY 22 20  0 */ (n175 & 1'b0) | ((n175 | 1'b0) & n181);
assign n69  = /* CARRY  7 20  3 */ (1'b0 & n39) | ((1'b0 | n39) & n68);
assign n138 = /* CARRY 16 12  2 */ (n99 & io_0_11_0) | ((n99 | io_0_11_0) & n137);
assign n254 = /* CARRY 21 20  3 */ (1'b0 & n172) | ((1'b0 | n172) & n232);
assign n255 = /* CARRY 22 20  2 */ (1'b0 & n173) | ((1'b0 | n173) & n230);
assign n71  = /* CARRY  7 20  5 */ (n41 & 1'b0) | ((n41 | 1'b0) & n70);
assign n136 = /* CARRY 16 12  0 */ (io_0_11_0 & n97) | ((io_0_11_0 | n97) & n128);
assign n256 = /* CARRY 21 20  1 */ (n162 & 1'b0) | ((n162 | 1'b0) & n233);
assign n257 = /* CARRY 18 11  4 */ (1'b0 & n112) | ((1'b0 | n112) & n240);
assign n142 = /* CARRY 16 12  6 */ (n103 & io_0_11_0) | ((n103 | io_0_11_0) & n141);
assign n176 = /* CARRY 21 20  7 */ (1'b0 & n164) | ((1'b0 | n164) & n234);
/* FF 18 11  6 */ assign n258 = n259;
/* FF 16 12  4 */ always @(posedge n4) if (n121) n101 <= n1 ? 1'b1 : n260;
/* FF 21 20  5 */ assign n261 = n262;
/* FF  7 21  2 */ assign n44 = n263;
/* FF 17 11  1 */ assign n114 = n264;
/* FF  7 19  2 */ assign n37 = n265;
/* FF 18 11  0 */ assign n266 = n267;
/* FF 24 22  5 */ always @(posedge io_0_27_1) if (1'b1) n86 <= 1'b0 ? 1'b0 : n269;
/* FF 16 14  5 */ assign n88 = n270;
/* FF 18 12  0 */ assign n271 = n272;
/* FF 18 11  2 */ assign n273 = n274;
/* FF 24 22  7 */ assign n22 = n275;
/* FF 18 12  2 */ assign n276 = n277;
/* FF  9 25  6 */ assign n33 = n278;
/* FF 16 14  1 */ assign n279 = n280;
/* FF 18 12  4 */ assign n281 = n282;
/* FF 16 11  3 */ always @(posedge n4) if (n121) n92 <= n1 ? 1'b1 : n283;
/* FF 21 21  0 */ assign n155 = n284;
/* FF 16 14  3 */ always @(posedge io_16_33_1) if (1'b1) n107 <= n108 ? 1'b0 : n285;
/* FF 18 12  6 */ assign n286 = n287;
/* FF 26 20  6 */ assign n165 = n288;
/* FF 16 11  1 */ assign n289 = n290;
/* FF 22 21  6 */ assign n174 = n291;
/* FF 24 25  5 */ assign n61 = n292;
/* FF 16 11  7 */ always @(posedge n4) if (n121) n96 <= n1 ? 1'b1 : n293;
/* FF 23 20  2 */ assign n59 = n294;
/* FF 22 21  4 */ assign n153 = n295;
/* FF 24 25  7 */ assign n65 = n296;
/* FF 19 12  5 */ assign n157 = n297;
/* FF 16 11  5 */ always @(posedge n4) if (n121) n94 <= n1 ? 1'b1 : n298;
/* FF 23 20  4 */ assign n66 = n299;
/* FF 18 10  7 */ assign n152 = n300;
/* FF 21 19  3 */ assign n301 = n302;
/* FF 24 21  4 */ assign n189 = n303;
/* FF  9 19  1 */ assign n63 = n304;
/* FF 23 20  6 */ assign n172 = n305;
/* FF 15 15  5 */ always @(posedge io_16_33_1) if (1'b1) n90 <= 1'b0 ? 1'b0 : n306;
/* FF  7 23  5 */ assign n48 = n307;
/* FF 22 21  0 */ assign n177 = n308;
/* FF 17 12  7 */ assign n135 = n309;
/* FF 18 10  5 */ assign n151 = n310;
/* FF 21 19  1 */ assign n311 = n312;
/* FF 17 12  5 */ assign n133 = n313;
/* FF 22 19  0 */ assign n314 = n315;
/* FF 22 22  6 */ assign n178 = n317;
/* FF 21 19  7 */ assign n318 = n319;
/* FF 17 12  3 */ assign n121 = n320;
/* FF 22 19  2 */ assign n321 = n322;
/* FF 20 19  7 */ assign n161 = n323;
/* FF 24 21  2 */ assign n179 = n324;
/* FF 21 19  5 */ assign n325 = n326;
/* FF 23 21  1 */ assign n184 = n327;
/* FF  1 23  0 */ assign n18 = n328;
/* FF 17 12  1 */ assign n130 = n329;
/* FF 22 19  4 */ assign n330 = n331;
/* FF 20 19  5 */ assign n159 = n332;
/* FF 22 20  5 */ assign n333 = n334;
/* FF 26 21  2 */ assign n190 = n335;
/* FF 22 18  7 */ assign n169 = n336;
/* FF 22 19  6 */ assign n337 = n338;
/* FF 22 20  7 */ assign n339 = n340;
/* FF  7 20  0 */ assign n341 = n342;
/* FF 22 18  5 */ assign n168 = n344;
/* FF 18 13  0 */ assign n154 = n345;
/* FF 22 20  1 */ assign n346 = n347;
/* FF 17 10  3 */ assign n112 = n348;
/* FF  7 20  2 */ always @(posedge n4) if (n18) n38 <= 1'b0 ? 1'b0 : n349;
/* FF 24 26  1 */ assign n192 = n350;
/* FF 16 20  4 */ always @(posedge io_0_27_1) if (1'b1) n58 <= 1'b0 ? 1'b0 : n351;
/* FF 16 12  3 */ always @(posedge n4) if (n121) n100 <= n1 ? 1'b1 : n352;
/* FF 11 24  7 */ assign io_0_11_0 = n353;
/* FF 22 20  3 */ assign n354 = n355;
/* FF 16 15  3 */ always @(posedge io_16_33_1) if (n109) n110 <= n108 ? 1'b0 : n356;
/* FF  6 21  2 */ assign n31 = n357;
/* FF  7 20  4 */ always @(posedge n4) if (n18) n40 <= 1'b0 ? 1'b0 : n358;
/* FF 21 20  2 */ assign n359 = n360;
/* FF 16 12  1 */ always @(posedge n4) if (n121) n98 <= n1 ? 1'b1 : n361;
/* FF 17 11  6 */ assign n1 = n362;
/* FF  7 21  7 */ always @(posedge n4) if (1'b1) io_0_18_0 <= 1'b0 ? 1'b0 : n363;
/* FF 24 20  1 */ assign n52 = n364;
/* FF  7 20  6 */ always @(posedge n4) if (n18) n42 <= 1'b0 ? 1'b0 : n365;
/* FF 21 20  0 */ assign n366 = n367;
/* FF 16 12  7 */ always @(posedge n4) if (n121) n104 <= n1 ? 1'b1 : n368;
/* FF 17 11  4 */ assign n117 = n369;
/* FF  7 21  5 */ always @(posedge n4) if (1'b1) io_0_17_0 <= 1'b0 ? 1'b0 : n370;
/* FF 21 20  6 */ assign n371 = n372;
/* FF 17 13  0 */ assign n143 = n373;
/* FF 18 11  5 */ assign n374 = n375;
/* FF 16 12  5 */ always @(posedge n4) if (n121) n102 <= n1 ? 1'b1 : n376;
/* FF 17 11  2 */ assign n115 = n377;
/* FF 21 20  4 */ assign n378 = n379;
/* FF  9 23  3 */ assign n30 = n380;
/* FF  7 19  3 */ always @(posedge n4) if (1'b1) io_0_17_1 <= 1'b0 ? 1'b0 : n381;
/* FF 26 19  7 */ assign n208 = n382;
/* FF 18 11  7 */ assign n383 = n384;
/* FF 17 11  0 */ assign n113 = n385;
/* FF  7 21  1 */ always @(posedge n4) if (1'b1) io_0_20_1 <= 1'b0 ? 1'b0 : n386;
/* FF  7 22  1 */ always @(posedge n4) if (1'b1) io_0_22_1 <= 1'b0 ? 1'b0 : n387;
/* FF 18 12  1 */ assign n388 = n389;
/* FF 24 17  5 */ assign n25 = n390;
/* FF 18 11  1 */ assign n391 = n392;
/* FF 16 14  4 */ assign n108 = n393;
/* FF 20 20  2 */ assign n162 = n394;
/* FF 18 12  3 */ assign n395 = n396;
/* FF 24 17  7 */ assign n75 = n397;
/* FF 18 11  3 */ assign n398 = n399;
/* FF  7 22  5 */ always @(posedge n4) if (1'b1) io_0_22_0 <= 1'b0 ? 1'b0 : n400;
/* FF 18 12  5 */ assign n401 = n402;
/* FF 16 11  2 */ always @(posedge n4) if (n121) n91 <= n1 ? 1'b1 : n403;
/* FF 16 14  0 */ assign n404 = n405;
/* FF  6 20  1 */ always @(posedge n4) if (n18) n27 <= 1'b0 ? 1'b0 : n407;
/* FF 18 12  7 */ assign n408 = n409;
/* FF 16 11  0 */ assign n410 = n411;
/* FF 21 18  3 */ assign n163 = n413;
/* FF 16 14  2 */ always @(posedge io_16_33_1) if (1'b1) n106 <= n108 ? 1'b0 : n414;
/* FF 16 11  6 */ always @(posedge n4) if (n121) n95 <= n1 ? 1'b1 : n415;
/* FF 18 10  2 */ assign n150 = n416;
/* FF 16 11  4 */ always @(posedge n4) if (n121) n93 <= n1 ? 1'b1 : n417;
/* FF 22 21  5 */ assign n175 = n418;
/* FF  7 23  0 */ assign n46 = n419;
/* FF 18 10  0 */ assign n149 = n420;
/* FF 18 23  7 */ always @(posedge io_0_27_1) if (1'b1) n80 <= 1'b0 ? 1'b0 : n421;
/* FF 22 21  3 */ assign n173 = n422;
/* FF  9 19  2 */ assign n85 = n423;
/* FF 17 12  6 */ assign n134 = n424;
/* FF  7 25  0 */ assign n50 = n425;
/* FF 23 21  6 */ assign n185 = n426;
/* FF 16 13  5 */ always @(posedge io_16_33_1) if (n88) n4 <= 1'b0 ? 1'b0 : n427;
/* FF  9 19  0 */ assign n62 = n428;
/* FF 21 19  2 */ assign n429 = n430;
/* FF 15 15  4 */ always @(posedge io_16_33_1) if (1'b1) n89 <= 1'b0 ? 1'b0 : n431;
/* FF 17 12  4 */ assign n132 = n432;
/* FF 18 10  4 */ always @(posedge n4) if (n150) n105 <= n1 ? 1'b1 : n433;
/* FF 24 21  7 */ assign n21 = n434;
/* FF 21 19  0 */ assign n435 = n436;
/* FF  7 23  6 */ assign n49 = n438;
/* FF 17 12  2 */ assign n131 = n439;
/* FF 22 19  1 */ assign n440 = n441;
/* FF 20 19  6 */ assign n160 = n442;
/* FF 21 19  6 */ assign n443 = n444;
/* FF 17 12  0 */ assign n129 = n445;
/* FF 22 19  3 */ assign n446 = n447;
/* FF 17 21  4 */ assign n120 = n448;
/* FF 23 21  0 */ assign n183 = n449;
/* FF 21 19  4 */ assign n450 = n451;
/* FF 24 21  3 */ assign n164 = n452;
/* FF 22 19  5 */ assign n453 = n454;
/* FF 22 20  4 */ assign n455 = n456;
/* FF 22 19  7 */ assign n457 = n458;
/* FF 22 20  6 */ assign n459 = n460;
/* FF 17 10  2 */ assign n111 = n461;
/* FF  7 20  1 */ assign n462 = n463;
/* FF 22 20  0 */ assign n464 = n465;
/* FF 16 15  2 */ assign n109 = n466;
/* FF  7 20  3 */ always @(posedge n4) if (n18) n39 <= 1'b0 ? 1'b0 : n467;
/* FF 30  1  6 */ assign io_31_0_1 = n468;
/* FF 24 26  0 */ assign n191 = n469;
/* FF 17 13  5 */ assign n145 = n470;
/* FF 22 18  2 */ assign n167 = n471;
/* FF 16 12  2 */ always @(posedge n4) if (n121) n99 <= n1 ? 1'b1 : n472;
/* FF 17 11  7 */ always @(posedge n4) if (n121) n119 <= n1 ? 1'b1 : n473;
/* FF 21 20  3 */ assign n474 = n475;
/* FF 22 20  2 */ assign n476 = n477;
/* FF  6 21  3 */ always @(posedge n4) if (n31) n32 <= 1'b0 ? 1'b0 : n478;
/* FF  7 20  5 */ always @(posedge n4) if (n18) n41 <= 1'b0 ? 1'b0 : n479;
/* FF 17 13  7 */ assign n146 = n480;
/* FF  7 19  4 */ assign n36 = n481;
/* FF 22 18  0 */ assign n166 = n482;
/* FF 16 12  0 */ always @(posedge n4) if (n121) n97 <= n1 ? 1'b1 : n483;
/* FF 12 23  0 */ assign io_0_16_0 = n484;
/* FF  7 21  6 */ assign n45 = n485;
/* FF 17 11  5 */ assign n118 = n486;
/* FF  7 20  7 */ always @(posedge n4) if (n18) n43 <= 1'b0 ? 1'b0 : n487;
/* FF 21 20  1 */ assign n488 = n489;
/* FF 18 11  4 */ assign n490 = n491;
/* FF 16 12  6 */ always @(posedge n4) if (n121) n103 <= n1 ? 1'b1 : n492;
/* FF 17 11  3 */ assign n116 = n493;
/* FF  7 21  4 */ always @(posedge n4) if (1'b1) io_0_20_0 <= 1'b0 ? 1'b0 : n494;
/* FF 21 20  7 */ assign n495 = n496;
/* FF 24 20  6 */ assign n171 = n497;
/* FF 17 13  3 */ assign n144 = n498;
/* FF  7 19  0 */ always @(posedge n4) if (1'b1) io_0_18_1 <= 1'b0 ? 1'b0 : n499;

endmodule

